// 
// Copyright 2015 Jeff Bush
// 
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
// 
//     http://www.apache.org/licenses/LICENSE-2.0
// 
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
// 

module gpio_controller
	#(parameter NUM_PINS = 8)

	(input				  clk,
	input				  reset,
	                      
	// IO bus interface   
	input [31:0]		  io_address,
	input				  io_read_en,	
	input [31:0]		  io_write_data,
	input				  io_write_en,
	output reg[31:0] 	  io_read_data,

	// To/from SD card
	inout[NUM_PINS - 1:0] gpio_value);	
	
	logic[NUM_PINS - 1:0] direction;
	logic[NUM_PINS - 1:0] output_value;

	genvar pin_idx;
	generate
	begin
		for (pin_idx = 0; pin_idx < NUM_PINS; pin_idx++)
		begin : pin_dir_gen
			assign gpio_value[pin_idx] = direction[pin_idx] 
				? output_value[pin_idx] : 1'bZ;
		end
	end
	
	synchronizer #(.WIDTH(NUM_PINS)) input_synchronizer(
		.data_o(io_read_data),
		.data_i(gpio_value),
		.*);
	
	always_ff @(posedge reset, posedge clk)
	begin
		if (reset)
		begin
			direction <= 0;
			output_value <= 0;
		end
		else if (io_write_en)
		begin
			if (io_address == 'h58)
				direction <= io_write_data;
			else if (io_address == 'h5c)
				output_value <= io_write_data;
		end
	end
endmodule
