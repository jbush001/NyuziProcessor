// 
// Copyright (C) 2011-2014 Jeff Bush
// 
// This library is free software; you can redistribute it and/or
// modify it under the terms of the GNU Library General Public
// License as published by the Free Software Foundation; either
// version 2 of the License, or (at your option) any later version.
// 
// This library is distributed in the hope that it will be useful,
// but WITHOUT ANY WARRANTY; without even the implied warranty of
// MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the GNU
// Library General Public License for more details.
// 
// You should have received a copy of the GNU Library General Public
// License along with this library; if not, write to the
// Free Software Foundation, Inc., 51 Franklin St, Fifth Floor,
// Boston, MA  02110-1301, USA.
// 


//
// This file is autogenerated by make_reciprocal_rom.py
//

module reciprocal_rom(
	input [5:0]        addr_i,
	output logic [5:0]   data_o);

	always_comb
	begin
		unique case (addr_i)
			6'h0: data_o = 6'h0;
			6'h1: data_o = 6'h3e;
			6'h2: data_o = 6'h3c;
			6'h3: data_o = 6'h3a;
			6'h4: data_o = 6'h38;
			6'h5: data_o = 6'h36;
			6'h6: data_o = 6'h35;
			6'h7: data_o = 6'h33;
			6'h8: data_o = 6'h31;
			6'h9: data_o = 6'h30;
			6'ha: data_o = 6'h2e;
			6'hb: data_o = 6'h2d;
			6'hc: data_o = 6'h2b;
			6'hd: data_o = 6'h2a;
			6'he: data_o = 6'h29;
			6'hf: data_o = 6'h27;
			6'h10: data_o = 6'h26;
			6'h11: data_o = 6'h25;
			6'h12: data_o = 6'h23;
			6'h13: data_o = 6'h22;
			6'h14: data_o = 6'h21;
			6'h15: data_o = 6'h20;
			6'h16: data_o = 6'h1f;
			6'h17: data_o = 6'h1e;
			6'h18: data_o = 6'h1d;
			6'h19: data_o = 6'h1c;
			6'h1a: data_o = 6'h1b;
			6'h1b: data_o = 6'h1a;
			6'h1c: data_o = 6'h19;
			6'h1d: data_o = 6'h18;
			6'h1e: data_o = 6'h17;
			6'h1f: data_o = 6'h16;
			6'h20: data_o = 6'h15;
			6'h21: data_o = 6'h14;
			6'h22: data_o = 6'h13;
			6'h23: data_o = 6'h12;
			6'h24: data_o = 6'h11;
			6'h25: data_o = 6'h11;
			6'h26: data_o = 6'h10;
			6'h27: data_o = 6'hf;
			6'h28: data_o = 6'he;
			6'h29: data_o = 6'he;
			6'h2a: data_o = 6'hd;
			6'h2b: data_o = 6'hc;
			6'h2c: data_o = 6'hb;
			6'h2d: data_o = 6'hb;
			6'h2e: data_o = 6'ha;
			6'h2f: data_o = 6'h9;
			6'h30: data_o = 6'h9;
			6'h31: data_o = 6'h8;
			6'h32: data_o = 6'h7;
			6'h33: data_o = 6'h7;
			6'h34: data_o = 6'h6;
			6'h35: data_o = 6'h6;
			6'h36: data_o = 6'h5;
			6'h37: data_o = 6'h4;
			6'h38: data_o = 6'h4;
			6'h39: data_o = 6'h3;
			6'h3a: data_o = 6'h3;
			6'h3b: data_o = 6'h2;
			6'h3c: data_o = 6'h2;
			6'h3d: data_o = 6'h1;
			6'h3e: data_o = 6'h1;
			6'h3f: data_o = 6'h0;
		endcase
	end
endmodule

// Local Variables:
// verilog-typedef-regexp:"_t$"
// End:

