// 
// Copyright 2011-2012 Jeff Bush
// 
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
// 
//     http://www.apache.org/licenses/LICENSE-2.0
// 
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
// 


//
// This file is autogenerated by make_reciprocal_rom.py
//

module reciprocal_rom(
	input [9:0]			addr_i,
	output reg [9:0]	data_o);

	always @*
	begin
		case (addr_i)
			10'h0: data_o = 10'h0; // 1.0 / 1.0 = 2.0
			10'h1: data_o = 10'h3fe; // 1.0 / 1.0009765625 = 1.998046875
			10'h2: data_o = 10'h3fc; // 1.0 / 1.001953125 = 1.99609375
			10'h3: data_o = 10'h3fa; // 1.0 / 1.0029296875 = 1.994140625
			10'h4: data_o = 10'h3f8; // 1.0 / 1.00390625 = 1.9921875
			10'h5: data_o = 10'h3f6; // 1.0 / 1.0048828125 = 1.990234375
			10'h6: data_o = 10'h3f4; // 1.0 / 1.005859375 = 1.98828125
			10'h7: data_o = 10'h3f2; // 1.0 / 1.0068359375 = 1.986328125
			10'h8: data_o = 10'h3f0; // 1.0 / 1.0078125 = 1.984375
			10'h9: data_o = 10'h3ee; // 1.0 / 1.0087890625 = 1.982421875
			10'ha: data_o = 10'h3ec; // 1.0 / 1.009765625 = 1.98046875
			10'hb: data_o = 10'h3ea; // 1.0 / 1.0107421875 = 1.978515625
			10'hc: data_o = 10'h3e8; // 1.0 / 1.01171875 = 1.9765625
			10'hd: data_o = 10'h3e6; // 1.0 / 1.0126953125 = 1.974609375
			10'he: data_o = 10'h3e4; // 1.0 / 1.013671875 = 1.97265625
			10'hf: data_o = 10'h3e2; // 1.0 / 1.0146484375 = 1.970703125
			10'h10: data_o = 10'h3e0; // 1.0 / 1.015625 = 1.96875
			10'h11: data_o = 10'h3de; // 1.0 / 1.0166015625 = 1.966796875
			10'h12: data_o = 10'h3dc; // 1.0 / 1.017578125 = 1.96484375
			10'h13: data_o = 10'h3da; // 1.0 / 1.0185546875 = 1.962890625
			10'h14: data_o = 10'h3d8; // 1.0 / 1.01953125 = 1.9609375
			10'h15: data_o = 10'h3d6; // 1.0 / 1.0205078125 = 1.958984375
			10'h16: data_o = 10'h3d4; // 1.0 / 1.021484375 = 1.95703125
			10'h17: data_o = 10'h3d3; // 1.0 / 1.0224609375 = 1.9560546875
			10'h18: data_o = 10'h3d1; // 1.0 / 1.0234375 = 1.9541015625
			10'h19: data_o = 10'h3cf; // 1.0 / 1.0244140625 = 1.9521484375
			10'h1a: data_o = 10'h3cd; // 1.0 / 1.025390625 = 1.9501953125
			10'h1b: data_o = 10'h3cb; // 1.0 / 1.0263671875 = 1.9482421875
			10'h1c: data_o = 10'h3c9; // 1.0 / 1.02734375 = 1.9462890625
			10'h1d: data_o = 10'h3c7; // 1.0 / 1.0283203125 = 1.9443359375
			10'h1e: data_o = 10'h3c5; // 1.0 / 1.029296875 = 1.9423828125
			10'h1f: data_o = 10'h3c3; // 1.0 / 1.0302734375 = 1.9404296875
			10'h20: data_o = 10'h3c1; // 1.0 / 1.03125 = 1.9384765625
			10'h21: data_o = 10'h3c0; // 1.0 / 1.0322265625 = 1.9375
			10'h22: data_o = 10'h3be; // 1.0 / 1.033203125 = 1.935546875
			10'h23: data_o = 10'h3bc; // 1.0 / 1.0341796875 = 1.93359375
			10'h24: data_o = 10'h3ba; // 1.0 / 1.03515625 = 1.931640625
			10'h25: data_o = 10'h3b8; // 1.0 / 1.0361328125 = 1.9296875
			10'h26: data_o = 10'h3b6; // 1.0 / 1.037109375 = 1.927734375
			10'h27: data_o = 10'h3b4; // 1.0 / 1.0380859375 = 1.92578125
			10'h28: data_o = 10'h3b3; // 1.0 / 1.0390625 = 1.9248046875
			10'h29: data_o = 10'h3b1; // 1.0 / 1.0400390625 = 1.9228515625
			10'h2a: data_o = 10'h3af; // 1.0 / 1.041015625 = 1.9208984375
			10'h2b: data_o = 10'h3ad; // 1.0 / 1.0419921875 = 1.9189453125
			10'h2c: data_o = 10'h3ab; // 1.0 / 1.04296875 = 1.9169921875
			10'h2d: data_o = 10'h3a9; // 1.0 / 1.0439453125 = 1.9150390625
			10'h2e: data_o = 10'h3a7; // 1.0 / 1.044921875 = 1.9130859375
			10'h2f: data_o = 10'h3a6; // 1.0 / 1.0458984375 = 1.912109375
			10'h30: data_o = 10'h3a4; // 1.0 / 1.046875 = 1.91015625
			10'h31: data_o = 10'h3a2; // 1.0 / 1.0478515625 = 1.908203125
			10'h32: data_o = 10'h3a0; // 1.0 / 1.048828125 = 1.90625
			10'h33: data_o = 10'h39e; // 1.0 / 1.0498046875 = 1.904296875
			10'h34: data_o = 10'h39d; // 1.0 / 1.05078125 = 1.9033203125
			10'h35: data_o = 10'h39b; // 1.0 / 1.0517578125 = 1.9013671875
			10'h36: data_o = 10'h399; // 1.0 / 1.052734375 = 1.8994140625
			10'h37: data_o = 10'h397; // 1.0 / 1.0537109375 = 1.8974609375
			10'h38: data_o = 10'h395; // 1.0 / 1.0546875 = 1.8955078125
			10'h39: data_o = 10'h394; // 1.0 / 1.0556640625 = 1.89453125
			10'h3a: data_o = 10'h392; // 1.0 / 1.056640625 = 1.892578125
			10'h3b: data_o = 10'h390; // 1.0 / 1.0576171875 = 1.890625
			10'h3c: data_o = 10'h38e; // 1.0 / 1.05859375 = 1.888671875
			10'h3d: data_o = 10'h38c; // 1.0 / 1.0595703125 = 1.88671875
			10'h3e: data_o = 10'h38b; // 1.0 / 1.060546875 = 1.8857421875
			10'h3f: data_o = 10'h389; // 1.0 / 1.0615234375 = 1.8837890625
			10'h40: data_o = 10'h387; // 1.0 / 1.0625 = 1.8818359375
			10'h41: data_o = 10'h385; // 1.0 / 1.0634765625 = 1.8798828125
			10'h42: data_o = 10'h383; // 1.0 / 1.064453125 = 1.8779296875
			10'h43: data_o = 10'h382; // 1.0 / 1.0654296875 = 1.876953125
			10'h44: data_o = 10'h380; // 1.0 / 1.06640625 = 1.875
			10'h45: data_o = 10'h37e; // 1.0 / 1.0673828125 = 1.873046875
			10'h46: data_o = 10'h37c; // 1.0 / 1.068359375 = 1.87109375
			10'h47: data_o = 10'h37b; // 1.0 / 1.0693359375 = 1.8701171875
			10'h48: data_o = 10'h379; // 1.0 / 1.0703125 = 1.8681640625
			10'h49: data_o = 10'h377; // 1.0 / 1.0712890625 = 1.8662109375
			10'h4a: data_o = 10'h375; // 1.0 / 1.072265625 = 1.8642578125
			10'h4b: data_o = 10'h374; // 1.0 / 1.0732421875 = 1.86328125
			10'h4c: data_o = 10'h372; // 1.0 / 1.07421875 = 1.861328125
			10'h4d: data_o = 10'h370; // 1.0 / 1.0751953125 = 1.859375
			10'h4e: data_o = 10'h36f; // 1.0 / 1.076171875 = 1.8583984375
			10'h4f: data_o = 10'h36d; // 1.0 / 1.0771484375 = 1.8564453125
			10'h50: data_o = 10'h36b; // 1.0 / 1.078125 = 1.8544921875
			10'h51: data_o = 10'h369; // 1.0 / 1.0791015625 = 1.8525390625
			10'h52: data_o = 10'h368; // 1.0 / 1.080078125 = 1.8515625
			10'h53: data_o = 10'h366; // 1.0 / 1.0810546875 = 1.849609375
			10'h54: data_o = 10'h364; // 1.0 / 1.08203125 = 1.84765625
			10'h55: data_o = 10'h363; // 1.0 / 1.0830078125 = 1.8466796875
			10'h56: data_o = 10'h361; // 1.0 / 1.083984375 = 1.8447265625
			10'h57: data_o = 10'h35f; // 1.0 / 1.0849609375 = 1.8427734375
			10'h58: data_o = 10'h35d; // 1.0 / 1.0859375 = 1.8408203125
			10'h59: data_o = 10'h35c; // 1.0 / 1.0869140625 = 1.83984375
			10'h5a: data_o = 10'h35a; // 1.0 / 1.087890625 = 1.837890625
			10'h5b: data_o = 10'h358; // 1.0 / 1.0888671875 = 1.8359375
			10'h5c: data_o = 10'h357; // 1.0 / 1.08984375 = 1.8349609375
			10'h5d: data_o = 10'h355; // 1.0 / 1.0908203125 = 1.8330078125
			10'h5e: data_o = 10'h353; // 1.0 / 1.091796875 = 1.8310546875
			10'h5f: data_o = 10'h352; // 1.0 / 1.0927734375 = 1.830078125
			10'h60: data_o = 10'h350; // 1.0 / 1.09375 = 1.828125
			10'h61: data_o = 10'h34e; // 1.0 / 1.0947265625 = 1.826171875
			10'h62: data_o = 10'h34d; // 1.0 / 1.095703125 = 1.8251953125
			10'h63: data_o = 10'h34b; // 1.0 / 1.0966796875 = 1.8232421875
			10'h64: data_o = 10'h349; // 1.0 / 1.09765625 = 1.8212890625
			10'h65: data_o = 10'h348; // 1.0 / 1.0986328125 = 1.8203125
			10'h66: data_o = 10'h346; // 1.0 / 1.099609375 = 1.818359375
			10'h67: data_o = 10'h344; // 1.0 / 1.1005859375 = 1.81640625
			10'h68: data_o = 10'h343; // 1.0 / 1.1015625 = 1.8154296875
			10'h69: data_o = 10'h341; // 1.0 / 1.1025390625 = 1.8134765625
			10'h6a: data_o = 10'h33f; // 1.0 / 1.103515625 = 1.8115234375
			10'h6b: data_o = 10'h33e; // 1.0 / 1.1044921875 = 1.810546875
			10'h6c: data_o = 10'h33c; // 1.0 / 1.10546875 = 1.80859375
			10'h6d: data_o = 10'h33a; // 1.0 / 1.1064453125 = 1.806640625
			10'h6e: data_o = 10'h339; // 1.0 / 1.107421875 = 1.8056640625
			10'h6f: data_o = 10'h337; // 1.0 / 1.1083984375 = 1.8037109375
			10'h70: data_o = 10'h336; // 1.0 / 1.109375 = 1.802734375
			10'h71: data_o = 10'h334; // 1.0 / 1.1103515625 = 1.80078125
			10'h72: data_o = 10'h332; // 1.0 / 1.111328125 = 1.798828125
			10'h73: data_o = 10'h331; // 1.0 / 1.1123046875 = 1.7978515625
			10'h74: data_o = 10'h32f; // 1.0 / 1.11328125 = 1.7958984375
			10'h75: data_o = 10'h32d; // 1.0 / 1.1142578125 = 1.7939453125
			10'h76: data_o = 10'h32c; // 1.0 / 1.115234375 = 1.79296875
			10'h77: data_o = 10'h32a; // 1.0 / 1.1162109375 = 1.791015625
			10'h78: data_o = 10'h329; // 1.0 / 1.1171875 = 1.7900390625
			10'h79: data_o = 10'h327; // 1.0 / 1.1181640625 = 1.7880859375
			10'h7a: data_o = 10'h325; // 1.0 / 1.119140625 = 1.7861328125
			10'h7b: data_o = 10'h324; // 1.0 / 1.1201171875 = 1.78515625
			10'h7c: data_o = 10'h322; // 1.0 / 1.12109375 = 1.783203125
			10'h7d: data_o = 10'h321; // 1.0 / 1.1220703125 = 1.7822265625
			10'h7e: data_o = 10'h31f; // 1.0 / 1.123046875 = 1.7802734375
			10'h7f: data_o = 10'h31e; // 1.0 / 1.1240234375 = 1.779296875
			10'h80: data_o = 10'h31c; // 1.0 / 1.125 = 1.77734375
			10'h81: data_o = 10'h31a; // 1.0 / 1.1259765625 = 1.775390625
			10'h82: data_o = 10'h319; // 1.0 / 1.126953125 = 1.7744140625
			10'h83: data_o = 10'h317; // 1.0 / 1.1279296875 = 1.7724609375
			10'h84: data_o = 10'h316; // 1.0 / 1.12890625 = 1.771484375
			10'h85: data_o = 10'h314; // 1.0 / 1.1298828125 = 1.76953125
			10'h86: data_o = 10'h313; // 1.0 / 1.130859375 = 1.7685546875
			10'h87: data_o = 10'h311; // 1.0 / 1.1318359375 = 1.7666015625
			10'h88: data_o = 10'h30f; // 1.0 / 1.1328125 = 1.7646484375
			10'h89: data_o = 10'h30e; // 1.0 / 1.1337890625 = 1.763671875
			10'h8a: data_o = 10'h30c; // 1.0 / 1.134765625 = 1.76171875
			10'h8b: data_o = 10'h30b; // 1.0 / 1.1357421875 = 1.7607421875
			10'h8c: data_o = 10'h309; // 1.0 / 1.13671875 = 1.7587890625
			10'h8d: data_o = 10'h308; // 1.0 / 1.1376953125 = 1.7578125
			10'h8e: data_o = 10'h306; // 1.0 / 1.138671875 = 1.755859375
			10'h8f: data_o = 10'h305; // 1.0 / 1.1396484375 = 1.7548828125
			10'h90: data_o = 10'h303; // 1.0 / 1.140625 = 1.7529296875
			10'h91: data_o = 10'h301; // 1.0 / 1.1416015625 = 1.7509765625
			10'h92: data_o = 10'h300; // 1.0 / 1.142578125 = 1.75
			10'h93: data_o = 10'h2fe; // 1.0 / 1.1435546875 = 1.748046875
			10'h94: data_o = 10'h2fd; // 1.0 / 1.14453125 = 1.7470703125
			10'h95: data_o = 10'h2fb; // 1.0 / 1.1455078125 = 1.7451171875
			10'h96: data_o = 10'h2fa; // 1.0 / 1.146484375 = 1.744140625
			10'h97: data_o = 10'h2f8; // 1.0 / 1.1474609375 = 1.7421875
			10'h98: data_o = 10'h2f7; // 1.0 / 1.1484375 = 1.7412109375
			10'h99: data_o = 10'h2f5; // 1.0 / 1.1494140625 = 1.7392578125
			10'h9a: data_o = 10'h2f4; // 1.0 / 1.150390625 = 1.73828125
			10'h9b: data_o = 10'h2f2; // 1.0 / 1.1513671875 = 1.736328125
			10'h9c: data_o = 10'h2f1; // 1.0 / 1.15234375 = 1.7353515625
			10'h9d: data_o = 10'h2ef; // 1.0 / 1.1533203125 = 1.7333984375
			10'h9e: data_o = 10'h2ee; // 1.0 / 1.154296875 = 1.732421875
			10'h9f: data_o = 10'h2ec; // 1.0 / 1.1552734375 = 1.73046875
			10'ha0: data_o = 10'h2eb; // 1.0 / 1.15625 = 1.7294921875
			10'ha1: data_o = 10'h2e9; // 1.0 / 1.1572265625 = 1.7275390625
			10'ha2: data_o = 10'h2e8; // 1.0 / 1.158203125 = 1.7265625
			10'ha3: data_o = 10'h2e6; // 1.0 / 1.1591796875 = 1.724609375
			10'ha4: data_o = 10'h2e5; // 1.0 / 1.16015625 = 1.7236328125
			10'ha5: data_o = 10'h2e3; // 1.0 / 1.1611328125 = 1.7216796875
			10'ha6: data_o = 10'h2e2; // 1.0 / 1.162109375 = 1.720703125
			10'ha7: data_o = 10'h2e0; // 1.0 / 1.1630859375 = 1.71875
			10'ha8: data_o = 10'h2df; // 1.0 / 1.1640625 = 1.7177734375
			10'ha9: data_o = 10'h2dd; // 1.0 / 1.1650390625 = 1.7158203125
			10'haa: data_o = 10'h2dc; // 1.0 / 1.166015625 = 1.71484375
			10'hab: data_o = 10'h2da; // 1.0 / 1.1669921875 = 1.712890625
			10'hac: data_o = 10'h2d9; // 1.0 / 1.16796875 = 1.7119140625
			10'had: data_o = 10'h2d8; // 1.0 / 1.1689453125 = 1.7109375
			10'hae: data_o = 10'h2d6; // 1.0 / 1.169921875 = 1.708984375
			10'haf: data_o = 10'h2d5; // 1.0 / 1.1708984375 = 1.7080078125
			10'hb0: data_o = 10'h2d3; // 1.0 / 1.171875 = 1.7060546875
			10'hb1: data_o = 10'h2d2; // 1.0 / 1.1728515625 = 1.705078125
			10'hb2: data_o = 10'h2d0; // 1.0 / 1.173828125 = 1.703125
			10'hb3: data_o = 10'h2cf; // 1.0 / 1.1748046875 = 1.7021484375
			10'hb4: data_o = 10'h2cd; // 1.0 / 1.17578125 = 1.7001953125
			10'hb5: data_o = 10'h2cc; // 1.0 / 1.1767578125 = 1.69921875
			10'hb6: data_o = 10'h2ca; // 1.0 / 1.177734375 = 1.697265625
			10'hb7: data_o = 10'h2c9; // 1.0 / 1.1787109375 = 1.6962890625
			10'hb8: data_o = 10'h2c8; // 1.0 / 1.1796875 = 1.6953125
			10'hb9: data_o = 10'h2c6; // 1.0 / 1.1806640625 = 1.693359375
			10'hba: data_o = 10'h2c5; // 1.0 / 1.181640625 = 1.6923828125
			10'hbb: data_o = 10'h2c3; // 1.0 / 1.1826171875 = 1.6904296875
			10'hbc: data_o = 10'h2c2; // 1.0 / 1.18359375 = 1.689453125
			10'hbd: data_o = 10'h2c0; // 1.0 / 1.1845703125 = 1.6875
			10'hbe: data_o = 10'h2bf; // 1.0 / 1.185546875 = 1.6865234375
			10'hbf: data_o = 10'h2be; // 1.0 / 1.1865234375 = 1.685546875
			10'hc0: data_o = 10'h2bc; // 1.0 / 1.1875 = 1.68359375
			10'hc1: data_o = 10'h2bb; // 1.0 / 1.1884765625 = 1.6826171875
			10'hc2: data_o = 10'h2b9; // 1.0 / 1.189453125 = 1.6806640625
			10'hc3: data_o = 10'h2b8; // 1.0 / 1.1904296875 = 1.6796875
			10'hc4: data_o = 10'h2b6; // 1.0 / 1.19140625 = 1.677734375
			10'hc5: data_o = 10'h2b5; // 1.0 / 1.1923828125 = 1.6767578125
			10'hc6: data_o = 10'h2b4; // 1.0 / 1.193359375 = 1.67578125
			10'hc7: data_o = 10'h2b2; // 1.0 / 1.1943359375 = 1.673828125
			10'hc8: data_o = 10'h2b1; // 1.0 / 1.1953125 = 1.6728515625
			10'hc9: data_o = 10'h2af; // 1.0 / 1.1962890625 = 1.6708984375
			10'hca: data_o = 10'h2ae; // 1.0 / 1.197265625 = 1.669921875
			10'hcb: data_o = 10'h2ad; // 1.0 / 1.1982421875 = 1.6689453125
			10'hcc: data_o = 10'h2ab; // 1.0 / 1.19921875 = 1.6669921875
			10'hcd: data_o = 10'h2aa; // 1.0 / 1.2001953125 = 1.666015625
			10'hce: data_o = 10'h2a9; // 1.0 / 1.201171875 = 1.6650390625
			10'hcf: data_o = 10'h2a7; // 1.0 / 1.2021484375 = 1.6630859375
			10'hd0: data_o = 10'h2a6; // 1.0 / 1.203125 = 1.662109375
			10'hd1: data_o = 10'h2a4; // 1.0 / 1.2041015625 = 1.66015625
			10'hd2: data_o = 10'h2a3; // 1.0 / 1.205078125 = 1.6591796875
			10'hd3: data_o = 10'h2a2; // 1.0 / 1.2060546875 = 1.658203125
			10'hd4: data_o = 10'h2a0; // 1.0 / 1.20703125 = 1.65625
			10'hd5: data_o = 10'h29f; // 1.0 / 1.2080078125 = 1.6552734375
			10'hd6: data_o = 10'h29d; // 1.0 / 1.208984375 = 1.6533203125
			10'hd7: data_o = 10'h29c; // 1.0 / 1.2099609375 = 1.65234375
			10'hd8: data_o = 10'h29b; // 1.0 / 1.2109375 = 1.6513671875
			10'hd9: data_o = 10'h299; // 1.0 / 1.2119140625 = 1.6494140625
			10'hda: data_o = 10'h298; // 1.0 / 1.212890625 = 1.6484375
			10'hdb: data_o = 10'h297; // 1.0 / 1.2138671875 = 1.6474609375
			10'hdc: data_o = 10'h295; // 1.0 / 1.21484375 = 1.6455078125
			10'hdd: data_o = 10'h294; // 1.0 / 1.2158203125 = 1.64453125
			10'hde: data_o = 10'h293; // 1.0 / 1.216796875 = 1.6435546875
			10'hdf: data_o = 10'h291; // 1.0 / 1.2177734375 = 1.6416015625
			10'he0: data_o = 10'h290; // 1.0 / 1.21875 = 1.640625
			10'he1: data_o = 10'h28f; // 1.0 / 1.2197265625 = 1.6396484375
			10'he2: data_o = 10'h28d; // 1.0 / 1.220703125 = 1.6376953125
			10'he3: data_o = 10'h28c; // 1.0 / 1.2216796875 = 1.63671875
			10'he4: data_o = 10'h28b; // 1.0 / 1.22265625 = 1.6357421875
			10'he5: data_o = 10'h289; // 1.0 / 1.2236328125 = 1.6337890625
			10'he6: data_o = 10'h288; // 1.0 / 1.224609375 = 1.6328125
			10'he7: data_o = 10'h287; // 1.0 / 1.2255859375 = 1.6318359375
			10'he8: data_o = 10'h285; // 1.0 / 1.2265625 = 1.6298828125
			10'he9: data_o = 10'h284; // 1.0 / 1.2275390625 = 1.62890625
			10'hea: data_o = 10'h283; // 1.0 / 1.228515625 = 1.6279296875
			10'heb: data_o = 10'h281; // 1.0 / 1.2294921875 = 1.6259765625
			10'hec: data_o = 10'h280; // 1.0 / 1.23046875 = 1.625
			10'hed: data_o = 10'h27f; // 1.0 / 1.2314453125 = 1.6240234375
			10'hee: data_o = 10'h27d; // 1.0 / 1.232421875 = 1.6220703125
			10'hef: data_o = 10'h27c; // 1.0 / 1.2333984375 = 1.62109375
			10'hf0: data_o = 10'h27b; // 1.0 / 1.234375 = 1.6201171875
			10'hf1: data_o = 10'h279; // 1.0 / 1.2353515625 = 1.6181640625
			10'hf2: data_o = 10'h278; // 1.0 / 1.236328125 = 1.6171875
			10'hf3: data_o = 10'h277; // 1.0 / 1.2373046875 = 1.6162109375
			10'hf4: data_o = 10'h275; // 1.0 / 1.23828125 = 1.6142578125
			10'hf5: data_o = 10'h274; // 1.0 / 1.2392578125 = 1.61328125
			10'hf6: data_o = 10'h273; // 1.0 / 1.240234375 = 1.6123046875
			10'hf7: data_o = 10'h272; // 1.0 / 1.2412109375 = 1.611328125
			10'hf8: data_o = 10'h270; // 1.0 / 1.2421875 = 1.609375
			10'hf9: data_o = 10'h26f; // 1.0 / 1.2431640625 = 1.6083984375
			10'hfa: data_o = 10'h26e; // 1.0 / 1.244140625 = 1.607421875
			10'hfb: data_o = 10'h26c; // 1.0 / 1.2451171875 = 1.60546875
			10'hfc: data_o = 10'h26b; // 1.0 / 1.24609375 = 1.6044921875
			10'hfd: data_o = 10'h26a; // 1.0 / 1.2470703125 = 1.603515625
			10'hfe: data_o = 10'h268; // 1.0 / 1.248046875 = 1.6015625
			10'hff: data_o = 10'h267; // 1.0 / 1.2490234375 = 1.6005859375
			10'h100: data_o = 10'h266; // 1.0 / 1.25 = 1.599609375
			10'h101: data_o = 10'h265; // 1.0 / 1.2509765625 = 1.5986328125
			10'h102: data_o = 10'h263; // 1.0 / 1.251953125 = 1.5966796875
			10'h103: data_o = 10'h262; // 1.0 / 1.2529296875 = 1.595703125
			10'h104: data_o = 10'h261; // 1.0 / 1.25390625 = 1.5947265625
			10'h105: data_o = 10'h260; // 1.0 / 1.2548828125 = 1.59375
			10'h106: data_o = 10'h25e; // 1.0 / 1.255859375 = 1.591796875
			10'h107: data_o = 10'h25d; // 1.0 / 1.2568359375 = 1.5908203125
			10'h108: data_o = 10'h25c; // 1.0 / 1.2578125 = 1.58984375
			10'h109: data_o = 10'h25a; // 1.0 / 1.2587890625 = 1.587890625
			10'h10a: data_o = 10'h259; // 1.0 / 1.259765625 = 1.5869140625
			10'h10b: data_o = 10'h258; // 1.0 / 1.2607421875 = 1.5859375
			10'h10c: data_o = 10'h257; // 1.0 / 1.26171875 = 1.5849609375
			10'h10d: data_o = 10'h255; // 1.0 / 1.2626953125 = 1.5830078125
			10'h10e: data_o = 10'h254; // 1.0 / 1.263671875 = 1.58203125
			10'h10f: data_o = 10'h253; // 1.0 / 1.2646484375 = 1.5810546875
			10'h110: data_o = 10'h252; // 1.0 / 1.265625 = 1.580078125
			10'h111: data_o = 10'h250; // 1.0 / 1.2666015625 = 1.578125
			10'h112: data_o = 10'h24f; // 1.0 / 1.267578125 = 1.5771484375
			10'h113: data_o = 10'h24e; // 1.0 / 1.2685546875 = 1.576171875
			10'h114: data_o = 10'h24d; // 1.0 / 1.26953125 = 1.5751953125
			10'h115: data_o = 10'h24b; // 1.0 / 1.2705078125 = 1.5732421875
			10'h116: data_o = 10'h24a; // 1.0 / 1.271484375 = 1.572265625
			10'h117: data_o = 10'h249; // 1.0 / 1.2724609375 = 1.5712890625
			10'h118: data_o = 10'h248; // 1.0 / 1.2734375 = 1.5703125
			10'h119: data_o = 10'h247; // 1.0 / 1.2744140625 = 1.5693359375
			10'h11a: data_o = 10'h245; // 1.0 / 1.275390625 = 1.5673828125
			10'h11b: data_o = 10'h244; // 1.0 / 1.2763671875 = 1.56640625
			10'h11c: data_o = 10'h243; // 1.0 / 1.27734375 = 1.5654296875
			10'h11d: data_o = 10'h242; // 1.0 / 1.2783203125 = 1.564453125
			10'h11e: data_o = 10'h240; // 1.0 / 1.279296875 = 1.5625
			10'h11f: data_o = 10'h23f; // 1.0 / 1.2802734375 = 1.5615234375
			10'h120: data_o = 10'h23e; // 1.0 / 1.28125 = 1.560546875
			10'h121: data_o = 10'h23d; // 1.0 / 1.2822265625 = 1.5595703125
			10'h122: data_o = 10'h23c; // 1.0 / 1.283203125 = 1.55859375
			10'h123: data_o = 10'h23a; // 1.0 / 1.2841796875 = 1.556640625
			10'h124: data_o = 10'h239; // 1.0 / 1.28515625 = 1.5556640625
			10'h125: data_o = 10'h238; // 1.0 / 1.2861328125 = 1.5546875
			10'h126: data_o = 10'h237; // 1.0 / 1.287109375 = 1.5537109375
			10'h127: data_o = 10'h235; // 1.0 / 1.2880859375 = 1.5517578125
			10'h128: data_o = 10'h234; // 1.0 / 1.2890625 = 1.55078125
			10'h129: data_o = 10'h233; // 1.0 / 1.2900390625 = 1.5498046875
			10'h12a: data_o = 10'h232; // 1.0 / 1.291015625 = 1.548828125
			10'h12b: data_o = 10'h231; // 1.0 / 1.2919921875 = 1.5478515625
			10'h12c: data_o = 10'h22f; // 1.0 / 1.29296875 = 1.5458984375
			10'h12d: data_o = 10'h22e; // 1.0 / 1.2939453125 = 1.544921875
			10'h12e: data_o = 10'h22d; // 1.0 / 1.294921875 = 1.5439453125
			10'h12f: data_o = 10'h22c; // 1.0 / 1.2958984375 = 1.54296875
			10'h130: data_o = 10'h22b; // 1.0 / 1.296875 = 1.5419921875
			10'h131: data_o = 10'h229; // 1.0 / 1.2978515625 = 1.5400390625
			10'h132: data_o = 10'h228; // 1.0 / 1.298828125 = 1.5390625
			10'h133: data_o = 10'h227; // 1.0 / 1.2998046875 = 1.5380859375
			10'h134: data_o = 10'h226; // 1.0 / 1.30078125 = 1.537109375
			10'h135: data_o = 10'h225; // 1.0 / 1.3017578125 = 1.5361328125
			10'h136: data_o = 10'h224; // 1.0 / 1.302734375 = 1.53515625
			10'h137: data_o = 10'h222; // 1.0 / 1.3037109375 = 1.533203125
			10'h138: data_o = 10'h221; // 1.0 / 1.3046875 = 1.5322265625
			10'h139: data_o = 10'h220; // 1.0 / 1.3056640625 = 1.53125
			10'h13a: data_o = 10'h21f; // 1.0 / 1.306640625 = 1.5302734375
			10'h13b: data_o = 10'h21e; // 1.0 / 1.3076171875 = 1.529296875
			10'h13c: data_o = 10'h21d; // 1.0 / 1.30859375 = 1.5283203125
			10'h13d: data_o = 10'h21b; // 1.0 / 1.3095703125 = 1.5263671875
			10'h13e: data_o = 10'h21a; // 1.0 / 1.310546875 = 1.525390625
			10'h13f: data_o = 10'h219; // 1.0 / 1.3115234375 = 1.5244140625
			10'h140: data_o = 10'h218; // 1.0 / 1.3125 = 1.5234375
			10'h141: data_o = 10'h217; // 1.0 / 1.3134765625 = 1.5224609375
			10'h142: data_o = 10'h216; // 1.0 / 1.314453125 = 1.521484375
			10'h143: data_o = 10'h214; // 1.0 / 1.3154296875 = 1.51953125
			10'h144: data_o = 10'h213; // 1.0 / 1.31640625 = 1.5185546875
			10'h145: data_o = 10'h212; // 1.0 / 1.3173828125 = 1.517578125
			10'h146: data_o = 10'h211; // 1.0 / 1.318359375 = 1.5166015625
			10'h147: data_o = 10'h210; // 1.0 / 1.3193359375 = 1.515625
			10'h148: data_o = 10'h20f; // 1.0 / 1.3203125 = 1.5146484375
			10'h149: data_o = 10'h20e; // 1.0 / 1.3212890625 = 1.513671875
			10'h14a: data_o = 10'h20c; // 1.0 / 1.322265625 = 1.51171875
			10'h14b: data_o = 10'h20b; // 1.0 / 1.3232421875 = 1.5107421875
			10'h14c: data_o = 10'h20a; // 1.0 / 1.32421875 = 1.509765625
			10'h14d: data_o = 10'h209; // 1.0 / 1.3251953125 = 1.5087890625
			10'h14e: data_o = 10'h208; // 1.0 / 1.326171875 = 1.5078125
			10'h14f: data_o = 10'h207; // 1.0 / 1.3271484375 = 1.5068359375
			10'h150: data_o = 10'h206; // 1.0 / 1.328125 = 1.505859375
			10'h151: data_o = 10'h204; // 1.0 / 1.3291015625 = 1.50390625
			10'h152: data_o = 10'h203; // 1.0 / 1.330078125 = 1.5029296875
			10'h153: data_o = 10'h202; // 1.0 / 1.3310546875 = 1.501953125
			10'h154: data_o = 10'h201; // 1.0 / 1.33203125 = 1.5009765625
			10'h155: data_o = 10'h200; // 1.0 / 1.3330078125 = 1.5
			10'h156: data_o = 10'h1ff; // 1.0 / 1.333984375 = 1.4990234375
			10'h157: data_o = 10'h1fe; // 1.0 / 1.3349609375 = 1.498046875
			10'h158: data_o = 10'h1fd; // 1.0 / 1.3359375 = 1.4970703125
			10'h159: data_o = 10'h1fb; // 1.0 / 1.3369140625 = 1.4951171875
			10'h15a: data_o = 10'h1fa; // 1.0 / 1.337890625 = 1.494140625
			10'h15b: data_o = 10'h1f9; // 1.0 / 1.3388671875 = 1.4931640625
			10'h15c: data_o = 10'h1f8; // 1.0 / 1.33984375 = 1.4921875
			10'h15d: data_o = 10'h1f7; // 1.0 / 1.3408203125 = 1.4912109375
			10'h15e: data_o = 10'h1f6; // 1.0 / 1.341796875 = 1.490234375
			10'h15f: data_o = 10'h1f5; // 1.0 / 1.3427734375 = 1.4892578125
			10'h160: data_o = 10'h1f4; // 1.0 / 1.34375 = 1.48828125
			10'h161: data_o = 10'h1f2; // 1.0 / 1.3447265625 = 1.486328125
			10'h162: data_o = 10'h1f1; // 1.0 / 1.345703125 = 1.4853515625
			10'h163: data_o = 10'h1f0; // 1.0 / 1.3466796875 = 1.484375
			10'h164: data_o = 10'h1ef; // 1.0 / 1.34765625 = 1.4833984375
			10'h165: data_o = 10'h1ee; // 1.0 / 1.3486328125 = 1.482421875
			10'h166: data_o = 10'h1ed; // 1.0 / 1.349609375 = 1.4814453125
			10'h167: data_o = 10'h1ec; // 1.0 / 1.3505859375 = 1.48046875
			10'h168: data_o = 10'h1eb; // 1.0 / 1.3515625 = 1.4794921875
			10'h169: data_o = 10'h1ea; // 1.0 / 1.3525390625 = 1.478515625
			10'h16a: data_o = 10'h1e9; // 1.0 / 1.353515625 = 1.4775390625
			10'h16b: data_o = 10'h1e8; // 1.0 / 1.3544921875 = 1.4765625
			10'h16c: data_o = 10'h1e6; // 1.0 / 1.35546875 = 1.474609375
			10'h16d: data_o = 10'h1e5; // 1.0 / 1.3564453125 = 1.4736328125
			10'h16e: data_o = 10'h1e4; // 1.0 / 1.357421875 = 1.47265625
			10'h16f: data_o = 10'h1e3; // 1.0 / 1.3583984375 = 1.4716796875
			10'h170: data_o = 10'h1e2; // 1.0 / 1.359375 = 1.470703125
			10'h171: data_o = 10'h1e1; // 1.0 / 1.3603515625 = 1.4697265625
			10'h172: data_o = 10'h1e0; // 1.0 / 1.361328125 = 1.46875
			10'h173: data_o = 10'h1df; // 1.0 / 1.3623046875 = 1.4677734375
			10'h174: data_o = 10'h1de; // 1.0 / 1.36328125 = 1.466796875
			10'h175: data_o = 10'h1dd; // 1.0 / 1.3642578125 = 1.4658203125
			10'h176: data_o = 10'h1dc; // 1.0 / 1.365234375 = 1.46484375
			10'h177: data_o = 10'h1db; // 1.0 / 1.3662109375 = 1.4638671875
			10'h178: data_o = 10'h1d9; // 1.0 / 1.3671875 = 1.4619140625
			10'h179: data_o = 10'h1d8; // 1.0 / 1.3681640625 = 1.4609375
			10'h17a: data_o = 10'h1d7; // 1.0 / 1.369140625 = 1.4599609375
			10'h17b: data_o = 10'h1d6; // 1.0 / 1.3701171875 = 1.458984375
			10'h17c: data_o = 10'h1d5; // 1.0 / 1.37109375 = 1.4580078125
			10'h17d: data_o = 10'h1d4; // 1.0 / 1.3720703125 = 1.45703125
			10'h17e: data_o = 10'h1d3; // 1.0 / 1.373046875 = 1.4560546875
			10'h17f: data_o = 10'h1d2; // 1.0 / 1.3740234375 = 1.455078125
			10'h180: data_o = 10'h1d1; // 1.0 / 1.375 = 1.4541015625
			10'h181: data_o = 10'h1d0; // 1.0 / 1.3759765625 = 1.453125
			10'h182: data_o = 10'h1cf; // 1.0 / 1.376953125 = 1.4521484375
			10'h183: data_o = 10'h1ce; // 1.0 / 1.3779296875 = 1.451171875
			10'h184: data_o = 10'h1cd; // 1.0 / 1.37890625 = 1.4501953125
			10'h185: data_o = 10'h1cc; // 1.0 / 1.3798828125 = 1.44921875
			10'h186: data_o = 10'h1cb; // 1.0 / 1.380859375 = 1.4482421875
			10'h187: data_o = 10'h1ca; // 1.0 / 1.3818359375 = 1.447265625
			10'h188: data_o = 10'h1c9; // 1.0 / 1.3828125 = 1.4462890625
			10'h189: data_o = 10'h1c7; // 1.0 / 1.3837890625 = 1.4443359375
			10'h18a: data_o = 10'h1c6; // 1.0 / 1.384765625 = 1.443359375
			10'h18b: data_o = 10'h1c5; // 1.0 / 1.3857421875 = 1.4423828125
			10'h18c: data_o = 10'h1c4; // 1.0 / 1.38671875 = 1.44140625
			10'h18d: data_o = 10'h1c3; // 1.0 / 1.3876953125 = 1.4404296875
			10'h18e: data_o = 10'h1c2; // 1.0 / 1.388671875 = 1.439453125
			10'h18f: data_o = 10'h1c1; // 1.0 / 1.3896484375 = 1.4384765625
			10'h190: data_o = 10'h1c0; // 1.0 / 1.390625 = 1.4375
			10'h191: data_o = 10'h1bf; // 1.0 / 1.3916015625 = 1.4365234375
			10'h192: data_o = 10'h1be; // 1.0 / 1.392578125 = 1.435546875
			10'h193: data_o = 10'h1bd; // 1.0 / 1.3935546875 = 1.4345703125
			10'h194: data_o = 10'h1bc; // 1.0 / 1.39453125 = 1.43359375
			10'h195: data_o = 10'h1bb; // 1.0 / 1.3955078125 = 1.4326171875
			10'h196: data_o = 10'h1ba; // 1.0 / 1.396484375 = 1.431640625
			10'h197: data_o = 10'h1b9; // 1.0 / 1.3974609375 = 1.4306640625
			10'h198: data_o = 10'h1b8; // 1.0 / 1.3984375 = 1.4296875
			10'h199: data_o = 10'h1b7; // 1.0 / 1.3994140625 = 1.4287109375
			10'h19a: data_o = 10'h1b6; // 1.0 / 1.400390625 = 1.427734375
			10'h19b: data_o = 10'h1b5; // 1.0 / 1.4013671875 = 1.4267578125
			10'h19c: data_o = 10'h1b4; // 1.0 / 1.40234375 = 1.42578125
			10'h19d: data_o = 10'h1b3; // 1.0 / 1.4033203125 = 1.4248046875
			10'h19e: data_o = 10'h1b2; // 1.0 / 1.404296875 = 1.423828125
			10'h19f: data_o = 10'h1b1; // 1.0 / 1.4052734375 = 1.4228515625
			10'h1a0: data_o = 10'h1b0; // 1.0 / 1.40625 = 1.421875
			10'h1a1: data_o = 10'h1af; // 1.0 / 1.4072265625 = 1.4208984375
			10'h1a2: data_o = 10'h1ae; // 1.0 / 1.408203125 = 1.419921875
			10'h1a3: data_o = 10'h1ad; // 1.0 / 1.4091796875 = 1.4189453125
			10'h1a4: data_o = 10'h1ac; // 1.0 / 1.41015625 = 1.41796875
			10'h1a5: data_o = 10'h1ab; // 1.0 / 1.4111328125 = 1.4169921875
			10'h1a6: data_o = 10'h1aa; // 1.0 / 1.412109375 = 1.416015625
			10'h1a7: data_o = 10'h1a9; // 1.0 / 1.4130859375 = 1.4150390625
			10'h1a8: data_o = 10'h1a8; // 1.0 / 1.4140625 = 1.4140625
			10'h1a9: data_o = 10'h1a7; // 1.0 / 1.4150390625 = 1.4130859375
			10'h1aa: data_o = 10'h1a6; // 1.0 / 1.416015625 = 1.412109375
			10'h1ab: data_o = 10'h1a5; // 1.0 / 1.4169921875 = 1.4111328125
			10'h1ac: data_o = 10'h1a4; // 1.0 / 1.41796875 = 1.41015625
			10'h1ad: data_o = 10'h1a3; // 1.0 / 1.4189453125 = 1.4091796875
			10'h1ae: data_o = 10'h1a2; // 1.0 / 1.419921875 = 1.408203125
			10'h1af: data_o = 10'h1a1; // 1.0 / 1.4208984375 = 1.4072265625
			10'h1b0: data_o = 10'h1a0; // 1.0 / 1.421875 = 1.40625
			10'h1b1: data_o = 10'h19f; // 1.0 / 1.4228515625 = 1.4052734375
			10'h1b2: data_o = 10'h19e; // 1.0 / 1.423828125 = 1.404296875
			10'h1b3: data_o = 10'h19d; // 1.0 / 1.4248046875 = 1.4033203125
			10'h1b4: data_o = 10'h19c; // 1.0 / 1.42578125 = 1.40234375
			10'h1b5: data_o = 10'h19b; // 1.0 / 1.4267578125 = 1.4013671875
			10'h1b6: data_o = 10'h19a; // 1.0 / 1.427734375 = 1.400390625
			10'h1b7: data_o = 10'h199; // 1.0 / 1.4287109375 = 1.3994140625
			10'h1b8: data_o = 10'h198; // 1.0 / 1.4296875 = 1.3984375
			10'h1b9: data_o = 10'h197; // 1.0 / 1.4306640625 = 1.3974609375
			10'h1ba: data_o = 10'h196; // 1.0 / 1.431640625 = 1.396484375
			10'h1bb: data_o = 10'h195; // 1.0 / 1.4326171875 = 1.3955078125
			10'h1bc: data_o = 10'h194; // 1.0 / 1.43359375 = 1.39453125
			10'h1bd: data_o = 10'h193; // 1.0 / 1.4345703125 = 1.3935546875
			10'h1be: data_o = 10'h192; // 1.0 / 1.435546875 = 1.392578125
			10'h1bf: data_o = 10'h191; // 1.0 / 1.4365234375 = 1.3916015625
			10'h1c0: data_o = 10'h190; // 1.0 / 1.4375 = 1.390625
			10'h1c1: data_o = 10'h18f; // 1.0 / 1.4384765625 = 1.3896484375
			10'h1c2: data_o = 10'h18e; // 1.0 / 1.439453125 = 1.388671875
			10'h1c3: data_o = 10'h18d; // 1.0 / 1.4404296875 = 1.3876953125
			10'h1c4: data_o = 10'h18c; // 1.0 / 1.44140625 = 1.38671875
			10'h1c5: data_o = 10'h18b; // 1.0 / 1.4423828125 = 1.3857421875
			10'h1c6: data_o = 10'h18a; // 1.0 / 1.443359375 = 1.384765625
			10'h1c7: data_o = 10'h189; // 1.0 / 1.4443359375 = 1.3837890625
			10'h1c8: data_o = 10'h188; // 1.0 / 1.4453125 = 1.3828125
			10'h1c9: data_o = 10'h188; // 1.0 / 1.4462890625 = 1.3828125
			10'h1ca: data_o = 10'h187; // 1.0 / 1.447265625 = 1.3818359375
			10'h1cb: data_o = 10'h186; // 1.0 / 1.4482421875 = 1.380859375
			10'h1cc: data_o = 10'h185; // 1.0 / 1.44921875 = 1.3798828125
			10'h1cd: data_o = 10'h184; // 1.0 / 1.4501953125 = 1.37890625
			10'h1ce: data_o = 10'h183; // 1.0 / 1.451171875 = 1.3779296875
			10'h1cf: data_o = 10'h182; // 1.0 / 1.4521484375 = 1.376953125
			10'h1d0: data_o = 10'h181; // 1.0 / 1.453125 = 1.3759765625
			10'h1d1: data_o = 10'h180; // 1.0 / 1.4541015625 = 1.375
			10'h1d2: data_o = 10'h17f; // 1.0 / 1.455078125 = 1.3740234375
			10'h1d3: data_o = 10'h17e; // 1.0 / 1.4560546875 = 1.373046875
			10'h1d4: data_o = 10'h17d; // 1.0 / 1.45703125 = 1.3720703125
			10'h1d5: data_o = 10'h17c; // 1.0 / 1.4580078125 = 1.37109375
			10'h1d6: data_o = 10'h17b; // 1.0 / 1.458984375 = 1.3701171875
			10'h1d7: data_o = 10'h17a; // 1.0 / 1.4599609375 = 1.369140625
			10'h1d8: data_o = 10'h179; // 1.0 / 1.4609375 = 1.3681640625
			10'h1d9: data_o = 10'h178; // 1.0 / 1.4619140625 = 1.3671875
			10'h1da: data_o = 10'h177; // 1.0 / 1.462890625 = 1.3662109375
			10'h1db: data_o = 10'h177; // 1.0 / 1.4638671875 = 1.3662109375
			10'h1dc: data_o = 10'h176; // 1.0 / 1.46484375 = 1.365234375
			10'h1dd: data_o = 10'h175; // 1.0 / 1.4658203125 = 1.3642578125
			10'h1de: data_o = 10'h174; // 1.0 / 1.466796875 = 1.36328125
			10'h1df: data_o = 10'h173; // 1.0 / 1.4677734375 = 1.3623046875
			10'h1e0: data_o = 10'h172; // 1.0 / 1.46875 = 1.361328125
			10'h1e1: data_o = 10'h171; // 1.0 / 1.4697265625 = 1.3603515625
			10'h1e2: data_o = 10'h170; // 1.0 / 1.470703125 = 1.359375
			10'h1e3: data_o = 10'h16f; // 1.0 / 1.4716796875 = 1.3583984375
			10'h1e4: data_o = 10'h16e; // 1.0 / 1.47265625 = 1.357421875
			10'h1e5: data_o = 10'h16d; // 1.0 / 1.4736328125 = 1.3564453125
			10'h1e6: data_o = 10'h16c; // 1.0 / 1.474609375 = 1.35546875
			10'h1e7: data_o = 10'h16b; // 1.0 / 1.4755859375 = 1.3544921875
			10'h1e8: data_o = 10'h16b; // 1.0 / 1.4765625 = 1.3544921875
			10'h1e9: data_o = 10'h16a; // 1.0 / 1.4775390625 = 1.353515625
			10'h1ea: data_o = 10'h169; // 1.0 / 1.478515625 = 1.3525390625
			10'h1eb: data_o = 10'h168; // 1.0 / 1.4794921875 = 1.3515625
			10'h1ec: data_o = 10'h167; // 1.0 / 1.48046875 = 1.3505859375
			10'h1ed: data_o = 10'h166; // 1.0 / 1.4814453125 = 1.349609375
			10'h1ee: data_o = 10'h165; // 1.0 / 1.482421875 = 1.3486328125
			10'h1ef: data_o = 10'h164; // 1.0 / 1.4833984375 = 1.34765625
			10'h1f0: data_o = 10'h163; // 1.0 / 1.484375 = 1.3466796875
			10'h1f1: data_o = 10'h162; // 1.0 / 1.4853515625 = 1.345703125
			10'h1f2: data_o = 10'h161; // 1.0 / 1.486328125 = 1.3447265625
			10'h1f3: data_o = 10'h160; // 1.0 / 1.4873046875 = 1.34375
			10'h1f4: data_o = 10'h160; // 1.0 / 1.48828125 = 1.34375
			10'h1f5: data_o = 10'h15f; // 1.0 / 1.4892578125 = 1.3427734375
			10'h1f6: data_o = 10'h15e; // 1.0 / 1.490234375 = 1.341796875
			10'h1f7: data_o = 10'h15d; // 1.0 / 1.4912109375 = 1.3408203125
			10'h1f8: data_o = 10'h15c; // 1.0 / 1.4921875 = 1.33984375
			10'h1f9: data_o = 10'h15b; // 1.0 / 1.4931640625 = 1.3388671875
			10'h1fa: data_o = 10'h15a; // 1.0 / 1.494140625 = 1.337890625
			10'h1fb: data_o = 10'h159; // 1.0 / 1.4951171875 = 1.3369140625
			10'h1fc: data_o = 10'h158; // 1.0 / 1.49609375 = 1.3359375
			10'h1fd: data_o = 10'h158; // 1.0 / 1.4970703125 = 1.3359375
			10'h1fe: data_o = 10'h157; // 1.0 / 1.498046875 = 1.3349609375
			10'h1ff: data_o = 10'h156; // 1.0 / 1.4990234375 = 1.333984375
			10'h200: data_o = 10'h155; // 1.0 / 1.5 = 1.3330078125
			10'h201: data_o = 10'h154; // 1.0 / 1.5009765625 = 1.33203125
			10'h202: data_o = 10'h153; // 1.0 / 1.501953125 = 1.3310546875
			10'h203: data_o = 10'h152; // 1.0 / 1.5029296875 = 1.330078125
			10'h204: data_o = 10'h151; // 1.0 / 1.50390625 = 1.3291015625
			10'h205: data_o = 10'h150; // 1.0 / 1.5048828125 = 1.328125
			10'h206: data_o = 10'h150; // 1.0 / 1.505859375 = 1.328125
			10'h207: data_o = 10'h14f; // 1.0 / 1.5068359375 = 1.3271484375
			10'h208: data_o = 10'h14e; // 1.0 / 1.5078125 = 1.326171875
			10'h209: data_o = 10'h14d; // 1.0 / 1.5087890625 = 1.3251953125
			10'h20a: data_o = 10'h14c; // 1.0 / 1.509765625 = 1.32421875
			10'h20b: data_o = 10'h14b; // 1.0 / 1.5107421875 = 1.3232421875
			10'h20c: data_o = 10'h14a; // 1.0 / 1.51171875 = 1.322265625
			10'h20d: data_o = 10'h149; // 1.0 / 1.5126953125 = 1.3212890625
			10'h20e: data_o = 10'h149; // 1.0 / 1.513671875 = 1.3212890625
			10'h20f: data_o = 10'h148; // 1.0 / 1.5146484375 = 1.3203125
			10'h210: data_o = 10'h147; // 1.0 / 1.515625 = 1.3193359375
			10'h211: data_o = 10'h146; // 1.0 / 1.5166015625 = 1.318359375
			10'h212: data_o = 10'h145; // 1.0 / 1.517578125 = 1.3173828125
			10'h213: data_o = 10'h144; // 1.0 / 1.5185546875 = 1.31640625
			10'h214: data_o = 10'h143; // 1.0 / 1.51953125 = 1.3154296875
			10'h215: data_o = 10'h142; // 1.0 / 1.5205078125 = 1.314453125
			10'h216: data_o = 10'h142; // 1.0 / 1.521484375 = 1.314453125
			10'h217: data_o = 10'h141; // 1.0 / 1.5224609375 = 1.3134765625
			10'h218: data_o = 10'h140; // 1.0 / 1.5234375 = 1.3125
			10'h219: data_o = 10'h13f; // 1.0 / 1.5244140625 = 1.3115234375
			10'h21a: data_o = 10'h13e; // 1.0 / 1.525390625 = 1.310546875
			10'h21b: data_o = 10'h13d; // 1.0 / 1.5263671875 = 1.3095703125
			10'h21c: data_o = 10'h13c; // 1.0 / 1.52734375 = 1.30859375
			10'h21d: data_o = 10'h13c; // 1.0 / 1.5283203125 = 1.30859375
			10'h21e: data_o = 10'h13b; // 1.0 / 1.529296875 = 1.3076171875
			10'h21f: data_o = 10'h13a; // 1.0 / 1.5302734375 = 1.306640625
			10'h220: data_o = 10'h139; // 1.0 / 1.53125 = 1.3056640625
			10'h221: data_o = 10'h138; // 1.0 / 1.5322265625 = 1.3046875
			10'h222: data_o = 10'h137; // 1.0 / 1.533203125 = 1.3037109375
			10'h223: data_o = 10'h136; // 1.0 / 1.5341796875 = 1.302734375
			10'h224: data_o = 10'h136; // 1.0 / 1.53515625 = 1.302734375
			10'h225: data_o = 10'h135; // 1.0 / 1.5361328125 = 1.3017578125
			10'h226: data_o = 10'h134; // 1.0 / 1.537109375 = 1.30078125
			10'h227: data_o = 10'h133; // 1.0 / 1.5380859375 = 1.2998046875
			10'h228: data_o = 10'h132; // 1.0 / 1.5390625 = 1.298828125
			10'h229: data_o = 10'h131; // 1.0 / 1.5400390625 = 1.2978515625
			10'h22a: data_o = 10'h130; // 1.0 / 1.541015625 = 1.296875
			10'h22b: data_o = 10'h130; // 1.0 / 1.5419921875 = 1.296875
			10'h22c: data_o = 10'h12f; // 1.0 / 1.54296875 = 1.2958984375
			10'h22d: data_o = 10'h12e; // 1.0 / 1.5439453125 = 1.294921875
			10'h22e: data_o = 10'h12d; // 1.0 / 1.544921875 = 1.2939453125
			10'h22f: data_o = 10'h12c; // 1.0 / 1.5458984375 = 1.29296875
			10'h230: data_o = 10'h12b; // 1.0 / 1.546875 = 1.2919921875
			10'h231: data_o = 10'h12b; // 1.0 / 1.5478515625 = 1.2919921875
			10'h232: data_o = 10'h12a; // 1.0 / 1.548828125 = 1.291015625
			10'h233: data_o = 10'h129; // 1.0 / 1.5498046875 = 1.2900390625
			10'h234: data_o = 10'h128; // 1.0 / 1.55078125 = 1.2890625
			10'h235: data_o = 10'h127; // 1.0 / 1.5517578125 = 1.2880859375
			10'h236: data_o = 10'h126; // 1.0 / 1.552734375 = 1.287109375
			10'h237: data_o = 10'h126; // 1.0 / 1.5537109375 = 1.287109375
			10'h238: data_o = 10'h125; // 1.0 / 1.5546875 = 1.2861328125
			10'h239: data_o = 10'h124; // 1.0 / 1.5556640625 = 1.28515625
			10'h23a: data_o = 10'h123; // 1.0 / 1.556640625 = 1.2841796875
			10'h23b: data_o = 10'h122; // 1.0 / 1.5576171875 = 1.283203125
			10'h23c: data_o = 10'h122; // 1.0 / 1.55859375 = 1.283203125
			10'h23d: data_o = 10'h121; // 1.0 / 1.5595703125 = 1.2822265625
			10'h23e: data_o = 10'h120; // 1.0 / 1.560546875 = 1.28125
			10'h23f: data_o = 10'h11f; // 1.0 / 1.5615234375 = 1.2802734375
			10'h240: data_o = 10'h11e; // 1.0 / 1.5625 = 1.279296875
			10'h241: data_o = 10'h11d; // 1.0 / 1.5634765625 = 1.2783203125
			10'h242: data_o = 10'h11d; // 1.0 / 1.564453125 = 1.2783203125
			10'h243: data_o = 10'h11c; // 1.0 / 1.5654296875 = 1.27734375
			10'h244: data_o = 10'h11b; // 1.0 / 1.56640625 = 1.2763671875
			10'h245: data_o = 10'h11a; // 1.0 / 1.5673828125 = 1.275390625
			10'h246: data_o = 10'h119; // 1.0 / 1.568359375 = 1.2744140625
			10'h247: data_o = 10'h119; // 1.0 / 1.5693359375 = 1.2744140625
			10'h248: data_o = 10'h118; // 1.0 / 1.5703125 = 1.2734375
			10'h249: data_o = 10'h117; // 1.0 / 1.5712890625 = 1.2724609375
			10'h24a: data_o = 10'h116; // 1.0 / 1.572265625 = 1.271484375
			10'h24b: data_o = 10'h115; // 1.0 / 1.5732421875 = 1.2705078125
			10'h24c: data_o = 10'h114; // 1.0 / 1.57421875 = 1.26953125
			10'h24d: data_o = 10'h114; // 1.0 / 1.5751953125 = 1.26953125
			10'h24e: data_o = 10'h113; // 1.0 / 1.576171875 = 1.2685546875
			10'h24f: data_o = 10'h112; // 1.0 / 1.5771484375 = 1.267578125
			10'h250: data_o = 10'h111; // 1.0 / 1.578125 = 1.2666015625
			10'h251: data_o = 10'h110; // 1.0 / 1.5791015625 = 1.265625
			10'h252: data_o = 10'h110; // 1.0 / 1.580078125 = 1.265625
			10'h253: data_o = 10'h10f; // 1.0 / 1.5810546875 = 1.2646484375
			10'h254: data_o = 10'h10e; // 1.0 / 1.58203125 = 1.263671875
			10'h255: data_o = 10'h10d; // 1.0 / 1.5830078125 = 1.2626953125
			10'h256: data_o = 10'h10c; // 1.0 / 1.583984375 = 1.26171875
			10'h257: data_o = 10'h10c; // 1.0 / 1.5849609375 = 1.26171875
			10'h258: data_o = 10'h10b; // 1.0 / 1.5859375 = 1.2607421875
			10'h259: data_o = 10'h10a; // 1.0 / 1.5869140625 = 1.259765625
			10'h25a: data_o = 10'h109; // 1.0 / 1.587890625 = 1.2587890625
			10'h25b: data_o = 10'h108; // 1.0 / 1.5888671875 = 1.2578125
			10'h25c: data_o = 10'h108; // 1.0 / 1.58984375 = 1.2578125
			10'h25d: data_o = 10'h107; // 1.0 / 1.5908203125 = 1.2568359375
			10'h25e: data_o = 10'h106; // 1.0 / 1.591796875 = 1.255859375
			10'h25f: data_o = 10'h105; // 1.0 / 1.5927734375 = 1.2548828125
			10'h260: data_o = 10'h105; // 1.0 / 1.59375 = 1.2548828125
			10'h261: data_o = 10'h104; // 1.0 / 1.5947265625 = 1.25390625
			10'h262: data_o = 10'h103; // 1.0 / 1.595703125 = 1.2529296875
			10'h263: data_o = 10'h102; // 1.0 / 1.5966796875 = 1.251953125
			10'h264: data_o = 10'h101; // 1.0 / 1.59765625 = 1.2509765625
			10'h265: data_o = 10'h101; // 1.0 / 1.5986328125 = 1.2509765625
			10'h266: data_o = 10'h100; // 1.0 / 1.599609375 = 1.25
			10'h267: data_o = 10'hff; // 1.0 / 1.6005859375 = 1.2490234375
			10'h268: data_o = 10'hfe; // 1.0 / 1.6015625 = 1.248046875
			10'h269: data_o = 10'hfd; // 1.0 / 1.6025390625 = 1.2470703125
			10'h26a: data_o = 10'hfd; // 1.0 / 1.603515625 = 1.2470703125
			10'h26b: data_o = 10'hfc; // 1.0 / 1.6044921875 = 1.24609375
			10'h26c: data_o = 10'hfb; // 1.0 / 1.60546875 = 1.2451171875
			10'h26d: data_o = 10'hfa; // 1.0 / 1.6064453125 = 1.244140625
			10'h26e: data_o = 10'hfa; // 1.0 / 1.607421875 = 1.244140625
			10'h26f: data_o = 10'hf9; // 1.0 / 1.6083984375 = 1.2431640625
			10'h270: data_o = 10'hf8; // 1.0 / 1.609375 = 1.2421875
			10'h271: data_o = 10'hf7; // 1.0 / 1.6103515625 = 1.2412109375
			10'h272: data_o = 10'hf7; // 1.0 / 1.611328125 = 1.2412109375
			10'h273: data_o = 10'hf6; // 1.0 / 1.6123046875 = 1.240234375
			10'h274: data_o = 10'hf5; // 1.0 / 1.61328125 = 1.2392578125
			10'h275: data_o = 10'hf4; // 1.0 / 1.6142578125 = 1.23828125
			10'h276: data_o = 10'hf3; // 1.0 / 1.615234375 = 1.2373046875
			10'h277: data_o = 10'hf3; // 1.0 / 1.6162109375 = 1.2373046875
			10'h278: data_o = 10'hf2; // 1.0 / 1.6171875 = 1.236328125
			10'h279: data_o = 10'hf1; // 1.0 / 1.6181640625 = 1.2353515625
			10'h27a: data_o = 10'hf0; // 1.0 / 1.619140625 = 1.234375
			10'h27b: data_o = 10'hf0; // 1.0 / 1.6201171875 = 1.234375
			10'h27c: data_o = 10'hef; // 1.0 / 1.62109375 = 1.2333984375
			10'h27d: data_o = 10'hee; // 1.0 / 1.6220703125 = 1.232421875
			10'h27e: data_o = 10'hed; // 1.0 / 1.623046875 = 1.2314453125
			10'h27f: data_o = 10'hed; // 1.0 / 1.6240234375 = 1.2314453125
			10'h280: data_o = 10'hec; // 1.0 / 1.625 = 1.23046875
			10'h281: data_o = 10'heb; // 1.0 / 1.6259765625 = 1.2294921875
			10'h282: data_o = 10'hea; // 1.0 / 1.626953125 = 1.228515625
			10'h283: data_o = 10'hea; // 1.0 / 1.6279296875 = 1.228515625
			10'h284: data_o = 10'he9; // 1.0 / 1.62890625 = 1.2275390625
			10'h285: data_o = 10'he8; // 1.0 / 1.6298828125 = 1.2265625
			10'h286: data_o = 10'he7; // 1.0 / 1.630859375 = 1.2255859375
			10'h287: data_o = 10'he7; // 1.0 / 1.6318359375 = 1.2255859375
			10'h288: data_o = 10'he6; // 1.0 / 1.6328125 = 1.224609375
			10'h289: data_o = 10'he5; // 1.0 / 1.6337890625 = 1.2236328125
			10'h28a: data_o = 10'he4; // 1.0 / 1.634765625 = 1.22265625
			10'h28b: data_o = 10'he4; // 1.0 / 1.6357421875 = 1.22265625
			10'h28c: data_o = 10'he3; // 1.0 / 1.63671875 = 1.2216796875
			10'h28d: data_o = 10'he2; // 1.0 / 1.6376953125 = 1.220703125
			10'h28e: data_o = 10'he1; // 1.0 / 1.638671875 = 1.2197265625
			10'h28f: data_o = 10'he1; // 1.0 / 1.6396484375 = 1.2197265625
			10'h290: data_o = 10'he0; // 1.0 / 1.640625 = 1.21875
			10'h291: data_o = 10'hdf; // 1.0 / 1.6416015625 = 1.2177734375
			10'h292: data_o = 10'hde; // 1.0 / 1.642578125 = 1.216796875
			10'h293: data_o = 10'hde; // 1.0 / 1.6435546875 = 1.216796875
			10'h294: data_o = 10'hdd; // 1.0 / 1.64453125 = 1.2158203125
			10'h295: data_o = 10'hdc; // 1.0 / 1.6455078125 = 1.21484375
			10'h296: data_o = 10'hdb; // 1.0 / 1.646484375 = 1.2138671875
			10'h297: data_o = 10'hdb; // 1.0 / 1.6474609375 = 1.2138671875
			10'h298: data_o = 10'hda; // 1.0 / 1.6484375 = 1.212890625
			10'h299: data_o = 10'hd9; // 1.0 / 1.6494140625 = 1.2119140625
			10'h29a: data_o = 10'hd8; // 1.0 / 1.650390625 = 1.2109375
			10'h29b: data_o = 10'hd8; // 1.0 / 1.6513671875 = 1.2109375
			10'h29c: data_o = 10'hd7; // 1.0 / 1.65234375 = 1.2099609375
			10'h29d: data_o = 10'hd6; // 1.0 / 1.6533203125 = 1.208984375
			10'h29e: data_o = 10'hd5; // 1.0 / 1.654296875 = 1.2080078125
			10'h29f: data_o = 10'hd5; // 1.0 / 1.6552734375 = 1.2080078125
			10'h2a0: data_o = 10'hd4; // 1.0 / 1.65625 = 1.20703125
			10'h2a1: data_o = 10'hd3; // 1.0 / 1.6572265625 = 1.2060546875
			10'h2a2: data_o = 10'hd3; // 1.0 / 1.658203125 = 1.2060546875
			10'h2a3: data_o = 10'hd2; // 1.0 / 1.6591796875 = 1.205078125
			10'h2a4: data_o = 10'hd1; // 1.0 / 1.66015625 = 1.2041015625
			10'h2a5: data_o = 10'hd0; // 1.0 / 1.6611328125 = 1.203125
			10'h2a6: data_o = 10'hd0; // 1.0 / 1.662109375 = 1.203125
			10'h2a7: data_o = 10'hcf; // 1.0 / 1.6630859375 = 1.2021484375
			10'h2a8: data_o = 10'hce; // 1.0 / 1.6640625 = 1.201171875
			10'h2a9: data_o = 10'hce; // 1.0 / 1.6650390625 = 1.201171875
			10'h2aa: data_o = 10'hcd; // 1.0 / 1.666015625 = 1.2001953125
			10'h2ab: data_o = 10'hcc; // 1.0 / 1.6669921875 = 1.19921875
			10'h2ac: data_o = 10'hcb; // 1.0 / 1.66796875 = 1.1982421875
			10'h2ad: data_o = 10'hcb; // 1.0 / 1.6689453125 = 1.1982421875
			10'h2ae: data_o = 10'hca; // 1.0 / 1.669921875 = 1.197265625
			10'h2af: data_o = 10'hc9; // 1.0 / 1.6708984375 = 1.1962890625
			10'h2b0: data_o = 10'hc8; // 1.0 / 1.671875 = 1.1953125
			10'h2b1: data_o = 10'hc8; // 1.0 / 1.6728515625 = 1.1953125
			10'h2b2: data_o = 10'hc7; // 1.0 / 1.673828125 = 1.1943359375
			10'h2b3: data_o = 10'hc6; // 1.0 / 1.6748046875 = 1.193359375
			10'h2b4: data_o = 10'hc6; // 1.0 / 1.67578125 = 1.193359375
			10'h2b5: data_o = 10'hc5; // 1.0 / 1.6767578125 = 1.1923828125
			10'h2b6: data_o = 10'hc4; // 1.0 / 1.677734375 = 1.19140625
			10'h2b7: data_o = 10'hc3; // 1.0 / 1.6787109375 = 1.1904296875
			10'h2b8: data_o = 10'hc3; // 1.0 / 1.6796875 = 1.1904296875
			10'h2b9: data_o = 10'hc2; // 1.0 / 1.6806640625 = 1.189453125
			10'h2ba: data_o = 10'hc1; // 1.0 / 1.681640625 = 1.1884765625
			10'h2bb: data_o = 10'hc1; // 1.0 / 1.6826171875 = 1.1884765625
			10'h2bc: data_o = 10'hc0; // 1.0 / 1.68359375 = 1.1875
			10'h2bd: data_o = 10'hbf; // 1.0 / 1.6845703125 = 1.1865234375
			10'h2be: data_o = 10'hbf; // 1.0 / 1.685546875 = 1.1865234375
			10'h2bf: data_o = 10'hbe; // 1.0 / 1.6865234375 = 1.185546875
			10'h2c0: data_o = 10'hbd; // 1.0 / 1.6875 = 1.1845703125
			10'h2c1: data_o = 10'hbc; // 1.0 / 1.6884765625 = 1.18359375
			10'h2c2: data_o = 10'hbc; // 1.0 / 1.689453125 = 1.18359375
			10'h2c3: data_o = 10'hbb; // 1.0 / 1.6904296875 = 1.1826171875
			10'h2c4: data_o = 10'hba; // 1.0 / 1.69140625 = 1.181640625
			10'h2c5: data_o = 10'hba; // 1.0 / 1.6923828125 = 1.181640625
			10'h2c6: data_o = 10'hb9; // 1.0 / 1.693359375 = 1.1806640625
			10'h2c7: data_o = 10'hb8; // 1.0 / 1.6943359375 = 1.1796875
			10'h2c8: data_o = 10'hb8; // 1.0 / 1.6953125 = 1.1796875
			10'h2c9: data_o = 10'hb7; // 1.0 / 1.6962890625 = 1.1787109375
			10'h2ca: data_o = 10'hb6; // 1.0 / 1.697265625 = 1.177734375
			10'h2cb: data_o = 10'hb5; // 1.0 / 1.6982421875 = 1.1767578125
			10'h2cc: data_o = 10'hb5; // 1.0 / 1.69921875 = 1.1767578125
			10'h2cd: data_o = 10'hb4; // 1.0 / 1.7001953125 = 1.17578125
			10'h2ce: data_o = 10'hb3; // 1.0 / 1.701171875 = 1.1748046875
			10'h2cf: data_o = 10'hb3; // 1.0 / 1.7021484375 = 1.1748046875
			10'h2d0: data_o = 10'hb2; // 1.0 / 1.703125 = 1.173828125
			10'h2d1: data_o = 10'hb1; // 1.0 / 1.7041015625 = 1.1728515625
			10'h2d2: data_o = 10'hb1; // 1.0 / 1.705078125 = 1.1728515625
			10'h2d3: data_o = 10'hb0; // 1.0 / 1.7060546875 = 1.171875
			10'h2d4: data_o = 10'haf; // 1.0 / 1.70703125 = 1.1708984375
			10'h2d5: data_o = 10'haf; // 1.0 / 1.7080078125 = 1.1708984375
			10'h2d6: data_o = 10'hae; // 1.0 / 1.708984375 = 1.169921875
			10'h2d7: data_o = 10'had; // 1.0 / 1.7099609375 = 1.1689453125
			10'h2d8: data_o = 10'had; // 1.0 / 1.7109375 = 1.1689453125
			10'h2d9: data_o = 10'hac; // 1.0 / 1.7119140625 = 1.16796875
			10'h2da: data_o = 10'hab; // 1.0 / 1.712890625 = 1.1669921875
			10'h2db: data_o = 10'haa; // 1.0 / 1.7138671875 = 1.166015625
			10'h2dc: data_o = 10'haa; // 1.0 / 1.71484375 = 1.166015625
			10'h2dd: data_o = 10'ha9; // 1.0 / 1.7158203125 = 1.1650390625
			10'h2de: data_o = 10'ha8; // 1.0 / 1.716796875 = 1.1640625
			10'h2df: data_o = 10'ha8; // 1.0 / 1.7177734375 = 1.1640625
			10'h2e0: data_o = 10'ha7; // 1.0 / 1.71875 = 1.1630859375
			10'h2e1: data_o = 10'ha6; // 1.0 / 1.7197265625 = 1.162109375
			10'h2e2: data_o = 10'ha6; // 1.0 / 1.720703125 = 1.162109375
			10'h2e3: data_o = 10'ha5; // 1.0 / 1.7216796875 = 1.1611328125
			10'h2e4: data_o = 10'ha4; // 1.0 / 1.72265625 = 1.16015625
			10'h2e5: data_o = 10'ha4; // 1.0 / 1.7236328125 = 1.16015625
			10'h2e6: data_o = 10'ha3; // 1.0 / 1.724609375 = 1.1591796875
			10'h2e7: data_o = 10'ha2; // 1.0 / 1.7255859375 = 1.158203125
			10'h2e8: data_o = 10'ha2; // 1.0 / 1.7265625 = 1.158203125
			10'h2e9: data_o = 10'ha1; // 1.0 / 1.7275390625 = 1.1572265625
			10'h2ea: data_o = 10'ha0; // 1.0 / 1.728515625 = 1.15625
			10'h2eb: data_o = 10'ha0; // 1.0 / 1.7294921875 = 1.15625
			10'h2ec: data_o = 10'h9f; // 1.0 / 1.73046875 = 1.1552734375
			10'h2ed: data_o = 10'h9e; // 1.0 / 1.7314453125 = 1.154296875
			10'h2ee: data_o = 10'h9e; // 1.0 / 1.732421875 = 1.154296875
			10'h2ef: data_o = 10'h9d; // 1.0 / 1.7333984375 = 1.1533203125
			10'h2f0: data_o = 10'h9c; // 1.0 / 1.734375 = 1.15234375
			10'h2f1: data_o = 10'h9c; // 1.0 / 1.7353515625 = 1.15234375
			10'h2f2: data_o = 10'h9b; // 1.0 / 1.736328125 = 1.1513671875
			10'h2f3: data_o = 10'h9a; // 1.0 / 1.7373046875 = 1.150390625
			10'h2f4: data_o = 10'h9a; // 1.0 / 1.73828125 = 1.150390625
			10'h2f5: data_o = 10'h99; // 1.0 / 1.7392578125 = 1.1494140625
			10'h2f6: data_o = 10'h98; // 1.0 / 1.740234375 = 1.1484375
			10'h2f7: data_o = 10'h98; // 1.0 / 1.7412109375 = 1.1484375
			10'h2f8: data_o = 10'h97; // 1.0 / 1.7421875 = 1.1474609375
			10'h2f9: data_o = 10'h96; // 1.0 / 1.7431640625 = 1.146484375
			10'h2fa: data_o = 10'h96; // 1.0 / 1.744140625 = 1.146484375
			10'h2fb: data_o = 10'h95; // 1.0 / 1.7451171875 = 1.1455078125
			10'h2fc: data_o = 10'h94; // 1.0 / 1.74609375 = 1.14453125
			10'h2fd: data_o = 10'h94; // 1.0 / 1.7470703125 = 1.14453125
			10'h2fe: data_o = 10'h93; // 1.0 / 1.748046875 = 1.1435546875
			10'h2ff: data_o = 10'h92; // 1.0 / 1.7490234375 = 1.142578125
			10'h300: data_o = 10'h92; // 1.0 / 1.75 = 1.142578125
			10'h301: data_o = 10'h91; // 1.0 / 1.7509765625 = 1.1416015625
			10'h302: data_o = 10'h90; // 1.0 / 1.751953125 = 1.140625
			10'h303: data_o = 10'h90; // 1.0 / 1.7529296875 = 1.140625
			10'h304: data_o = 10'h8f; // 1.0 / 1.75390625 = 1.1396484375
			10'h305: data_o = 10'h8f; // 1.0 / 1.7548828125 = 1.1396484375
			10'h306: data_o = 10'h8e; // 1.0 / 1.755859375 = 1.138671875
			10'h307: data_o = 10'h8d; // 1.0 / 1.7568359375 = 1.1376953125
			10'h308: data_o = 10'h8d; // 1.0 / 1.7578125 = 1.1376953125
			10'h309: data_o = 10'h8c; // 1.0 / 1.7587890625 = 1.13671875
			10'h30a: data_o = 10'h8b; // 1.0 / 1.759765625 = 1.1357421875
			10'h30b: data_o = 10'h8b; // 1.0 / 1.7607421875 = 1.1357421875
			10'h30c: data_o = 10'h8a; // 1.0 / 1.76171875 = 1.134765625
			10'h30d: data_o = 10'h89; // 1.0 / 1.7626953125 = 1.1337890625
			10'h30e: data_o = 10'h89; // 1.0 / 1.763671875 = 1.1337890625
			10'h30f: data_o = 10'h88; // 1.0 / 1.7646484375 = 1.1328125
			10'h310: data_o = 10'h87; // 1.0 / 1.765625 = 1.1318359375
			10'h311: data_o = 10'h87; // 1.0 / 1.7666015625 = 1.1318359375
			10'h312: data_o = 10'h86; // 1.0 / 1.767578125 = 1.130859375
			10'h313: data_o = 10'h86; // 1.0 / 1.7685546875 = 1.130859375
			10'h314: data_o = 10'h85; // 1.0 / 1.76953125 = 1.1298828125
			10'h315: data_o = 10'h84; // 1.0 / 1.7705078125 = 1.12890625
			10'h316: data_o = 10'h84; // 1.0 / 1.771484375 = 1.12890625
			10'h317: data_o = 10'h83; // 1.0 / 1.7724609375 = 1.1279296875
			10'h318: data_o = 10'h82; // 1.0 / 1.7734375 = 1.126953125
			10'h319: data_o = 10'h82; // 1.0 / 1.7744140625 = 1.126953125
			10'h31a: data_o = 10'h81; // 1.0 / 1.775390625 = 1.1259765625
			10'h31b: data_o = 10'h80; // 1.0 / 1.7763671875 = 1.125
			10'h31c: data_o = 10'h80; // 1.0 / 1.77734375 = 1.125
			10'h31d: data_o = 10'h7f; // 1.0 / 1.7783203125 = 1.1240234375
			10'h31e: data_o = 10'h7f; // 1.0 / 1.779296875 = 1.1240234375
			10'h31f: data_o = 10'h7e; // 1.0 / 1.7802734375 = 1.123046875
			10'h320: data_o = 10'h7d; // 1.0 / 1.78125 = 1.1220703125
			10'h321: data_o = 10'h7d; // 1.0 / 1.7822265625 = 1.1220703125
			10'h322: data_o = 10'h7c; // 1.0 / 1.783203125 = 1.12109375
			10'h323: data_o = 10'h7b; // 1.0 / 1.7841796875 = 1.1201171875
			10'h324: data_o = 10'h7b; // 1.0 / 1.78515625 = 1.1201171875
			10'h325: data_o = 10'h7a; // 1.0 / 1.7861328125 = 1.119140625
			10'h326: data_o = 10'h79; // 1.0 / 1.787109375 = 1.1181640625
			10'h327: data_o = 10'h79; // 1.0 / 1.7880859375 = 1.1181640625
			10'h328: data_o = 10'h78; // 1.0 / 1.7890625 = 1.1171875
			10'h329: data_o = 10'h78; // 1.0 / 1.7900390625 = 1.1171875
			10'h32a: data_o = 10'h77; // 1.0 / 1.791015625 = 1.1162109375
			10'h32b: data_o = 10'h76; // 1.0 / 1.7919921875 = 1.115234375
			10'h32c: data_o = 10'h76; // 1.0 / 1.79296875 = 1.115234375
			10'h32d: data_o = 10'h75; // 1.0 / 1.7939453125 = 1.1142578125
			10'h32e: data_o = 10'h74; // 1.0 / 1.794921875 = 1.11328125
			10'h32f: data_o = 10'h74; // 1.0 / 1.7958984375 = 1.11328125
			10'h330: data_o = 10'h73; // 1.0 / 1.796875 = 1.1123046875
			10'h331: data_o = 10'h73; // 1.0 / 1.7978515625 = 1.1123046875
			10'h332: data_o = 10'h72; // 1.0 / 1.798828125 = 1.111328125
			10'h333: data_o = 10'h71; // 1.0 / 1.7998046875 = 1.1103515625
			10'h334: data_o = 10'h71; // 1.0 / 1.80078125 = 1.1103515625
			10'h335: data_o = 10'h70; // 1.0 / 1.8017578125 = 1.109375
			10'h336: data_o = 10'h70; // 1.0 / 1.802734375 = 1.109375
			10'h337: data_o = 10'h6f; // 1.0 / 1.8037109375 = 1.1083984375
			10'h338: data_o = 10'h6e; // 1.0 / 1.8046875 = 1.107421875
			10'h339: data_o = 10'h6e; // 1.0 / 1.8056640625 = 1.107421875
			10'h33a: data_o = 10'h6d; // 1.0 / 1.806640625 = 1.1064453125
			10'h33b: data_o = 10'h6c; // 1.0 / 1.8076171875 = 1.10546875
			10'h33c: data_o = 10'h6c; // 1.0 / 1.80859375 = 1.10546875
			10'h33d: data_o = 10'h6b; // 1.0 / 1.8095703125 = 1.1044921875
			10'h33e: data_o = 10'h6b; // 1.0 / 1.810546875 = 1.1044921875
			10'h33f: data_o = 10'h6a; // 1.0 / 1.8115234375 = 1.103515625
			10'h340: data_o = 10'h69; // 1.0 / 1.8125 = 1.1025390625
			10'h341: data_o = 10'h69; // 1.0 / 1.8134765625 = 1.1025390625
			10'h342: data_o = 10'h68; // 1.0 / 1.814453125 = 1.1015625
			10'h343: data_o = 10'h68; // 1.0 / 1.8154296875 = 1.1015625
			10'h344: data_o = 10'h67; // 1.0 / 1.81640625 = 1.1005859375
			10'h345: data_o = 10'h66; // 1.0 / 1.8173828125 = 1.099609375
			10'h346: data_o = 10'h66; // 1.0 / 1.818359375 = 1.099609375
			10'h347: data_o = 10'h65; // 1.0 / 1.8193359375 = 1.0986328125
			10'h348: data_o = 10'h65; // 1.0 / 1.8203125 = 1.0986328125
			10'h349: data_o = 10'h64; // 1.0 / 1.8212890625 = 1.09765625
			10'h34a: data_o = 10'h63; // 1.0 / 1.822265625 = 1.0966796875
			10'h34b: data_o = 10'h63; // 1.0 / 1.8232421875 = 1.0966796875
			10'h34c: data_o = 10'h62; // 1.0 / 1.82421875 = 1.095703125
			10'h34d: data_o = 10'h62; // 1.0 / 1.8251953125 = 1.095703125
			10'h34e: data_o = 10'h61; // 1.0 / 1.826171875 = 1.0947265625
			10'h34f: data_o = 10'h60; // 1.0 / 1.8271484375 = 1.09375
			10'h350: data_o = 10'h60; // 1.0 / 1.828125 = 1.09375
			10'h351: data_o = 10'h5f; // 1.0 / 1.8291015625 = 1.0927734375
			10'h352: data_o = 10'h5f; // 1.0 / 1.830078125 = 1.0927734375
			10'h353: data_o = 10'h5e; // 1.0 / 1.8310546875 = 1.091796875
			10'h354: data_o = 10'h5d; // 1.0 / 1.83203125 = 1.0908203125
			10'h355: data_o = 10'h5d; // 1.0 / 1.8330078125 = 1.0908203125
			10'h356: data_o = 10'h5c; // 1.0 / 1.833984375 = 1.08984375
			10'h357: data_o = 10'h5c; // 1.0 / 1.8349609375 = 1.08984375
			10'h358: data_o = 10'h5b; // 1.0 / 1.8359375 = 1.0888671875
			10'h359: data_o = 10'h5a; // 1.0 / 1.8369140625 = 1.087890625
			10'h35a: data_o = 10'h5a; // 1.0 / 1.837890625 = 1.087890625
			10'h35b: data_o = 10'h59; // 1.0 / 1.8388671875 = 1.0869140625
			10'h35c: data_o = 10'h59; // 1.0 / 1.83984375 = 1.0869140625
			10'h35d: data_o = 10'h58; // 1.0 / 1.8408203125 = 1.0859375
			10'h35e: data_o = 10'h57; // 1.0 / 1.841796875 = 1.0849609375
			10'h35f: data_o = 10'h57; // 1.0 / 1.8427734375 = 1.0849609375
			10'h360: data_o = 10'h56; // 1.0 / 1.84375 = 1.083984375
			10'h361: data_o = 10'h56; // 1.0 / 1.8447265625 = 1.083984375
			10'h362: data_o = 10'h55; // 1.0 / 1.845703125 = 1.0830078125
			10'h363: data_o = 10'h55; // 1.0 / 1.8466796875 = 1.0830078125
			10'h364: data_o = 10'h54; // 1.0 / 1.84765625 = 1.08203125
			10'h365: data_o = 10'h53; // 1.0 / 1.8486328125 = 1.0810546875
			10'h366: data_o = 10'h53; // 1.0 / 1.849609375 = 1.0810546875
			10'h367: data_o = 10'h52; // 1.0 / 1.8505859375 = 1.080078125
			10'h368: data_o = 10'h52; // 1.0 / 1.8515625 = 1.080078125
			10'h369: data_o = 10'h51; // 1.0 / 1.8525390625 = 1.0791015625
			10'h36a: data_o = 10'h50; // 1.0 / 1.853515625 = 1.078125
			10'h36b: data_o = 10'h50; // 1.0 / 1.8544921875 = 1.078125
			10'h36c: data_o = 10'h4f; // 1.0 / 1.85546875 = 1.0771484375
			10'h36d: data_o = 10'h4f; // 1.0 / 1.8564453125 = 1.0771484375
			10'h36e: data_o = 10'h4e; // 1.0 / 1.857421875 = 1.076171875
			10'h36f: data_o = 10'h4e; // 1.0 / 1.8583984375 = 1.076171875
			10'h370: data_o = 10'h4d; // 1.0 / 1.859375 = 1.0751953125
			10'h371: data_o = 10'h4c; // 1.0 / 1.8603515625 = 1.07421875
			10'h372: data_o = 10'h4c; // 1.0 / 1.861328125 = 1.07421875
			10'h373: data_o = 10'h4b; // 1.0 / 1.8623046875 = 1.0732421875
			10'h374: data_o = 10'h4b; // 1.0 / 1.86328125 = 1.0732421875
			10'h375: data_o = 10'h4a; // 1.0 / 1.8642578125 = 1.072265625
			10'h376: data_o = 10'h49; // 1.0 / 1.865234375 = 1.0712890625
			10'h377: data_o = 10'h49; // 1.0 / 1.8662109375 = 1.0712890625
			10'h378: data_o = 10'h48; // 1.0 / 1.8671875 = 1.0703125
			10'h379: data_o = 10'h48; // 1.0 / 1.8681640625 = 1.0703125
			10'h37a: data_o = 10'h47; // 1.0 / 1.869140625 = 1.0693359375
			10'h37b: data_o = 10'h47; // 1.0 / 1.8701171875 = 1.0693359375
			10'h37c: data_o = 10'h46; // 1.0 / 1.87109375 = 1.068359375
			10'h37d: data_o = 10'h45; // 1.0 / 1.8720703125 = 1.0673828125
			10'h37e: data_o = 10'h45; // 1.0 / 1.873046875 = 1.0673828125
			10'h37f: data_o = 10'h44; // 1.0 / 1.8740234375 = 1.06640625
			10'h380: data_o = 10'h44; // 1.0 / 1.875 = 1.06640625
			10'h381: data_o = 10'h43; // 1.0 / 1.8759765625 = 1.0654296875
			10'h382: data_o = 10'h43; // 1.0 / 1.876953125 = 1.0654296875
			10'h383: data_o = 10'h42; // 1.0 / 1.8779296875 = 1.064453125
			10'h384: data_o = 10'h41; // 1.0 / 1.87890625 = 1.0634765625
			10'h385: data_o = 10'h41; // 1.0 / 1.8798828125 = 1.0634765625
			10'h386: data_o = 10'h40; // 1.0 / 1.880859375 = 1.0625
			10'h387: data_o = 10'h40; // 1.0 / 1.8818359375 = 1.0625
			10'h388: data_o = 10'h3f; // 1.0 / 1.8828125 = 1.0615234375
			10'h389: data_o = 10'h3f; // 1.0 / 1.8837890625 = 1.0615234375
			10'h38a: data_o = 10'h3e; // 1.0 / 1.884765625 = 1.060546875
			10'h38b: data_o = 10'h3e; // 1.0 / 1.8857421875 = 1.060546875
			10'h38c: data_o = 10'h3d; // 1.0 / 1.88671875 = 1.0595703125
			10'h38d: data_o = 10'h3c; // 1.0 / 1.8876953125 = 1.05859375
			10'h38e: data_o = 10'h3c; // 1.0 / 1.888671875 = 1.05859375
			10'h38f: data_o = 10'h3b; // 1.0 / 1.8896484375 = 1.0576171875
			10'h390: data_o = 10'h3b; // 1.0 / 1.890625 = 1.0576171875
			10'h391: data_o = 10'h3a; // 1.0 / 1.8916015625 = 1.056640625
			10'h392: data_o = 10'h3a; // 1.0 / 1.892578125 = 1.056640625
			10'h393: data_o = 10'h39; // 1.0 / 1.8935546875 = 1.0556640625
			10'h394: data_o = 10'h39; // 1.0 / 1.89453125 = 1.0556640625
			10'h395: data_o = 10'h38; // 1.0 / 1.8955078125 = 1.0546875
			10'h396: data_o = 10'h37; // 1.0 / 1.896484375 = 1.0537109375
			10'h397: data_o = 10'h37; // 1.0 / 1.8974609375 = 1.0537109375
			10'h398: data_o = 10'h36; // 1.0 / 1.8984375 = 1.052734375
			10'h399: data_o = 10'h36; // 1.0 / 1.8994140625 = 1.052734375
			10'h39a: data_o = 10'h35; // 1.0 / 1.900390625 = 1.0517578125
			10'h39b: data_o = 10'h35; // 1.0 / 1.9013671875 = 1.0517578125
			10'h39c: data_o = 10'h34; // 1.0 / 1.90234375 = 1.05078125
			10'h39d: data_o = 10'h34; // 1.0 / 1.9033203125 = 1.05078125
			10'h39e: data_o = 10'h33; // 1.0 / 1.904296875 = 1.0498046875
			10'h39f: data_o = 10'h32; // 1.0 / 1.9052734375 = 1.048828125
			10'h3a0: data_o = 10'h32; // 1.0 / 1.90625 = 1.048828125
			10'h3a1: data_o = 10'h31; // 1.0 / 1.9072265625 = 1.0478515625
			10'h3a2: data_o = 10'h31; // 1.0 / 1.908203125 = 1.0478515625
			10'h3a3: data_o = 10'h30; // 1.0 / 1.9091796875 = 1.046875
			10'h3a4: data_o = 10'h30; // 1.0 / 1.91015625 = 1.046875
			10'h3a5: data_o = 10'h2f; // 1.0 / 1.9111328125 = 1.0458984375
			10'h3a6: data_o = 10'h2f; // 1.0 / 1.912109375 = 1.0458984375
			10'h3a7: data_o = 10'h2e; // 1.0 / 1.9130859375 = 1.044921875
			10'h3a8: data_o = 10'h2d; // 1.0 / 1.9140625 = 1.0439453125
			10'h3a9: data_o = 10'h2d; // 1.0 / 1.9150390625 = 1.0439453125
			10'h3aa: data_o = 10'h2c; // 1.0 / 1.916015625 = 1.04296875
			10'h3ab: data_o = 10'h2c; // 1.0 / 1.9169921875 = 1.04296875
			10'h3ac: data_o = 10'h2b; // 1.0 / 1.91796875 = 1.0419921875
			10'h3ad: data_o = 10'h2b; // 1.0 / 1.9189453125 = 1.0419921875
			10'h3ae: data_o = 10'h2a; // 1.0 / 1.919921875 = 1.041015625
			10'h3af: data_o = 10'h2a; // 1.0 / 1.9208984375 = 1.041015625
			10'h3b0: data_o = 10'h29; // 1.0 / 1.921875 = 1.0400390625
			10'h3b1: data_o = 10'h29; // 1.0 / 1.9228515625 = 1.0400390625
			10'h3b2: data_o = 10'h28; // 1.0 / 1.923828125 = 1.0390625
			10'h3b3: data_o = 10'h28; // 1.0 / 1.9248046875 = 1.0390625
			10'h3b4: data_o = 10'h27; // 1.0 / 1.92578125 = 1.0380859375
			10'h3b5: data_o = 10'h26; // 1.0 / 1.9267578125 = 1.037109375
			10'h3b6: data_o = 10'h26; // 1.0 / 1.927734375 = 1.037109375
			10'h3b7: data_o = 10'h25; // 1.0 / 1.9287109375 = 1.0361328125
			10'h3b8: data_o = 10'h25; // 1.0 / 1.9296875 = 1.0361328125
			10'h3b9: data_o = 10'h24; // 1.0 / 1.9306640625 = 1.03515625
			10'h3ba: data_o = 10'h24; // 1.0 / 1.931640625 = 1.03515625
			10'h3bb: data_o = 10'h23; // 1.0 / 1.9326171875 = 1.0341796875
			10'h3bc: data_o = 10'h23; // 1.0 / 1.93359375 = 1.0341796875
			10'h3bd: data_o = 10'h22; // 1.0 / 1.9345703125 = 1.033203125
			10'h3be: data_o = 10'h22; // 1.0 / 1.935546875 = 1.033203125
			10'h3bf: data_o = 10'h21; // 1.0 / 1.9365234375 = 1.0322265625
			10'h3c0: data_o = 10'h21; // 1.0 / 1.9375 = 1.0322265625
			10'h3c1: data_o = 10'h20; // 1.0 / 1.9384765625 = 1.03125
			10'h3c2: data_o = 10'h1f; // 1.0 / 1.939453125 = 1.0302734375
			10'h3c3: data_o = 10'h1f; // 1.0 / 1.9404296875 = 1.0302734375
			10'h3c4: data_o = 10'h1e; // 1.0 / 1.94140625 = 1.029296875
			10'h3c5: data_o = 10'h1e; // 1.0 / 1.9423828125 = 1.029296875
			10'h3c6: data_o = 10'h1d; // 1.0 / 1.943359375 = 1.0283203125
			10'h3c7: data_o = 10'h1d; // 1.0 / 1.9443359375 = 1.0283203125
			10'h3c8: data_o = 10'h1c; // 1.0 / 1.9453125 = 1.02734375
			10'h3c9: data_o = 10'h1c; // 1.0 / 1.9462890625 = 1.02734375
			10'h3ca: data_o = 10'h1b; // 1.0 / 1.947265625 = 1.0263671875
			10'h3cb: data_o = 10'h1b; // 1.0 / 1.9482421875 = 1.0263671875
			10'h3cc: data_o = 10'h1a; // 1.0 / 1.94921875 = 1.025390625
			10'h3cd: data_o = 10'h1a; // 1.0 / 1.9501953125 = 1.025390625
			10'h3ce: data_o = 10'h19; // 1.0 / 1.951171875 = 1.0244140625
			10'h3cf: data_o = 10'h19; // 1.0 / 1.9521484375 = 1.0244140625
			10'h3d0: data_o = 10'h18; // 1.0 / 1.953125 = 1.0234375
			10'h3d1: data_o = 10'h18; // 1.0 / 1.9541015625 = 1.0234375
			10'h3d2: data_o = 10'h17; // 1.0 / 1.955078125 = 1.0224609375
			10'h3d3: data_o = 10'h17; // 1.0 / 1.9560546875 = 1.0224609375
			10'h3d4: data_o = 10'h16; // 1.0 / 1.95703125 = 1.021484375
			10'h3d5: data_o = 10'h15; // 1.0 / 1.9580078125 = 1.0205078125
			10'h3d6: data_o = 10'h15; // 1.0 / 1.958984375 = 1.0205078125
			10'h3d7: data_o = 10'h14; // 1.0 / 1.9599609375 = 1.01953125
			10'h3d8: data_o = 10'h14; // 1.0 / 1.9609375 = 1.01953125
			10'h3d9: data_o = 10'h13; // 1.0 / 1.9619140625 = 1.0185546875
			10'h3da: data_o = 10'h13; // 1.0 / 1.962890625 = 1.0185546875
			10'h3db: data_o = 10'h12; // 1.0 / 1.9638671875 = 1.017578125
			10'h3dc: data_o = 10'h12; // 1.0 / 1.96484375 = 1.017578125
			10'h3dd: data_o = 10'h11; // 1.0 / 1.9658203125 = 1.0166015625
			10'h3de: data_o = 10'h11; // 1.0 / 1.966796875 = 1.0166015625
			10'h3df: data_o = 10'h10; // 1.0 / 1.9677734375 = 1.015625
			10'h3e0: data_o = 10'h10; // 1.0 / 1.96875 = 1.015625
			10'h3e1: data_o = 10'hf; // 1.0 / 1.9697265625 = 1.0146484375
			10'h3e2: data_o = 10'hf; // 1.0 / 1.970703125 = 1.0146484375
			10'h3e3: data_o = 10'he; // 1.0 / 1.9716796875 = 1.013671875
			10'h3e4: data_o = 10'he; // 1.0 / 1.97265625 = 1.013671875
			10'h3e5: data_o = 10'hd; // 1.0 / 1.9736328125 = 1.0126953125
			10'h3e6: data_o = 10'hd; // 1.0 / 1.974609375 = 1.0126953125
			10'h3e7: data_o = 10'hc; // 1.0 / 1.9755859375 = 1.01171875
			10'h3e8: data_o = 10'hc; // 1.0 / 1.9765625 = 1.01171875
			10'h3e9: data_o = 10'hb; // 1.0 / 1.9775390625 = 1.0107421875
			10'h3ea: data_o = 10'hb; // 1.0 / 1.978515625 = 1.0107421875
			10'h3eb: data_o = 10'ha; // 1.0 / 1.9794921875 = 1.009765625
			10'h3ec: data_o = 10'ha; // 1.0 / 1.98046875 = 1.009765625
			10'h3ed: data_o = 10'h9; // 1.0 / 1.9814453125 = 1.0087890625
			10'h3ee: data_o = 10'h9; // 1.0 / 1.982421875 = 1.0087890625
			10'h3ef: data_o = 10'h8; // 1.0 / 1.9833984375 = 1.0078125
			10'h3f0: data_o = 10'h8; // 1.0 / 1.984375 = 1.0078125
			10'h3f1: data_o = 10'h7; // 1.0 / 1.9853515625 = 1.0068359375
			10'h3f2: data_o = 10'h7; // 1.0 / 1.986328125 = 1.0068359375
			10'h3f3: data_o = 10'h6; // 1.0 / 1.9873046875 = 1.005859375
			10'h3f4: data_o = 10'h6; // 1.0 / 1.98828125 = 1.005859375
			10'h3f5: data_o = 10'h5; // 1.0 / 1.9892578125 = 1.0048828125
			10'h3f6: data_o = 10'h5; // 1.0 / 1.990234375 = 1.0048828125
			10'h3f7: data_o = 10'h4; // 1.0 / 1.9912109375 = 1.00390625
			10'h3f8: data_o = 10'h4; // 1.0 / 1.9921875 = 1.00390625
			10'h3f9: data_o = 10'h3; // 1.0 / 1.9931640625 = 1.0029296875
			10'h3fa: data_o = 10'h3; // 1.0 / 1.994140625 = 1.0029296875
			10'h3fb: data_o = 10'h2; // 1.0 / 1.9951171875 = 1.001953125
			10'h3fc: data_o = 10'h2; // 1.0 / 1.99609375 = 1.001953125
			10'h3fd: data_o = 10'h1; // 1.0 / 1.9970703125 = 1.0009765625
			10'h3fe: data_o = 10'h1; // 1.0 / 1.998046875 = 1.0009765625
			10'h3ff: data_o = 10'h0; // 1.0 / 1.9990234375 = 1.0
		endcase
	end
endmodule

