//
// Keep 4 instruction FIFOs (one for each strand) loaded.
//

module instruction_fetch_stage(
	input							clk,
	output reg[31:0]				icache_addr,
	input [31:0]					icache_data,
	input                           icache_hit,
	output							icache_request,
	output reg[1:0]					icache_req_strand = 0,
	input [3:0]						icache_load_complete_strands,
	input							icache_load_collision,

	output [31:0]					if_instruction0,
	output							if_instruction_valid0,
	output [31:0]					if_pc0,
	input							ss_instruction_req0,
	input							rb_rollback_strand0,
	input [31:0]					rb_rollback_pc0,

	output [31:0]					if_instruction1,
	output							if_instruction_valid1,
	output [31:0]					if_pc1,
	input							ss_instruction_req1,
	input							rb_rollback_strand1,
	input [31:0]					rb_rollback_pc1,

	output [31:0]					if_instruction2,
	output							if_instruction_valid2,
	output [31:0]					if_pc2,
	input							ss_instruction_req2,
	input							rb_rollback_strand2,
	input [31:0]					rb_rollback_pc2,

	output [31:0]					if_instruction3,
	output							if_instruction_valid3,
	output [31:0]					if_pc3,
	input							ss_instruction_req3,
	input							rb_rollback_strand3,
	input [31:0]					rb_rollback_pc3);
	
	reg[31:0]						program_counter0_ff = 0;
	reg[31:0]						program_counter0_nxt = 0;
	reg[31:0]						program_counter1_ff = 0;
	reg[31:0]						program_counter1_nxt = 0;
	reg[31:0]						program_counter2_ff = 0;
	reg[31:0]						program_counter2_nxt = 0;
	reg[31:0]						program_counter3_ff = 0;
	reg[31:0]						program_counter3_nxt = 0;
	wire							request0;
	wire							request1;
	wire							request2;
	wire							request3;
	reg[3:0]						instruction_cache_wait_ff = 0;
	reg[3:0]						instruction_cache_wait_nxt = 0;

	// This stores the last strand that issued a request to the cache (since results
	// have one cycle of latency, we need to remember this).
	reg[3:0]						cache_request_ff = 0;
	wire[3:0]						cache_request_nxt;

	// Issue least recently issued strand.  Don't issue strands that we know are
	// waiting on the cache.
	arbiter4 request_arb(
		.clk(clk),
		.req0_i(request0 & !instruction_cache_wait_nxt[0]),
		.req1_i(request1 & !instruction_cache_wait_nxt[1]),
		.req2_i(request2 & !instruction_cache_wait_nxt[2]),
		.req3_i(request3 & !instruction_cache_wait_nxt[3]),
		.update_lru_i(1'b1),
		.grant0_o(cache_request_nxt[0]),
		.grant1_o(cache_request_nxt[1]),
		.grant2_o(cache_request_nxt[2]),
		.grant3_o(cache_request_nxt[3]));
	
	assign icache_request = |cache_request_nxt;

	always @*
	begin
		case (cache_request_nxt)
			4'b1000: icache_addr = program_counter3_nxt;
			4'b0100: icache_addr = program_counter2_nxt;
			4'b0010: icache_addr = program_counter1_nxt;
			4'b0001: icache_addr = program_counter0_nxt;
			4'b0000: icache_addr = program_counter0_nxt;	// Don't care
			default: icache_addr = {32{1'bx}};	// Shouldn't happen
		endcase
	end

	always @*
	begin
		case (cache_request_nxt)
			4'b1000: icache_req_strand	 = 3;
			4'b0100: icache_req_strand	 = 2;
			4'b0010: icache_req_strand	 = 1;
			4'b0001: icache_req_strand	 = 0;
			4'b0000: icache_req_strand 	 = 0;	// Don't care
			default: icache_req_strand	 = {2{1'bx}};	// Shouldn't happen
		endcase
	end
	
	// Keep track of which strands are waiting on an icache fetch.
	always @*
	begin
		if (!icache_hit && cache_request_ff && !icache_load_collision)
		begin
			instruction_cache_wait_nxt = (instruction_cache_wait_ff & ~icache_load_complete_strands)
				| cache_request_ff;
		end
		else
		begin
			instruction_cache_wait_nxt = instruction_cache_wait_ff
				& ~icache_load_complete_strands;
		end
	end

	sync_fifo if0(
		.clk(clk),
		.flush_i(rb_rollback_strand0),
		.can_enqueue_o(request0),
		.enqueue_i(icache_hit && cache_request_ff[0]),
		.value_i({ program_counter0_nxt, icache_data[7:0], icache_data[15:8], 
			icache_data[23:16], icache_data[31:24] }),
		.can_dequeue_o(if_instruction_valid0),
		.dequeue_i(ss_instruction_req0 && if_instruction_valid0),	// FIXME instruction_valid_o is redundant
		.value_o({ if_pc0, if_instruction0 }));

	sync_fifo if1(
		.clk(clk),
		.flush_i(rb_rollback_strand1),
		.can_enqueue_o(request1),
		.enqueue_i(icache_hit && cache_request_ff[1]),
		.value_i({ program_counter1_nxt, icache_data[7:0], icache_data[15:8], 
			icache_data[23:16], icache_data[31:24] }),
		.can_dequeue_o(if_instruction_valid1),
		.dequeue_i(ss_instruction_req1 && if_instruction_valid1),	// FIXME instruction_valid_o is redundant
		.value_o({ if_pc1, if_instruction1 }));

	sync_fifo if2(
		.clk(clk),
		.flush_i(rb_rollback_strand2),
		.can_enqueue_o(request2),
		.enqueue_i(icache_hit && cache_request_ff[2]),
		.value_i({ program_counter2_nxt, icache_data[7:0], icache_data[15:8], 
			icache_data[23:16], icache_data[31:24] }),
		.can_dequeue_o(if_instruction_valid2),
		.dequeue_i(ss_instruction_req2 && if_instruction_valid2),	// FIXME instruction_valid_o is redundant
		.value_o({ if_pc2, if_instruction2 }));

	sync_fifo if3(
		.clk(clk),
		.flush_i(rb_rollback_strand3),
		.can_enqueue_o(request3),
		.enqueue_i(icache_hit && cache_request_ff[3]),
		.value_i({ program_counter3_nxt, icache_data[7:0], icache_data[15:8], 
			icache_data[23:16], icache_data[31:24] }),
		.can_dequeue_o(if_instruction_valid3),
		.dequeue_i(ss_instruction_req3 && if_instruction_valid3),	// FIXME instruction_valid_o is redundant
		.value_o({ if_pc3, if_instruction3 }));

	always @*
	begin
		if (rb_rollback_strand0)
			program_counter0_nxt = rb_rollback_pc0;
		else if (!icache_hit || !cache_request_ff[0])	
			program_counter0_nxt = program_counter0_ff;
		else
			program_counter0_nxt = program_counter0_ff + 32'd4;
	end

	always @*
	begin
		if (rb_rollback_strand1)
			program_counter1_nxt = rb_rollback_pc1;
		else if (!icache_hit || !cache_request_ff[1])	
			program_counter1_nxt = program_counter1_ff;
		else
			program_counter1_nxt = program_counter1_ff + 32'd4;
	end

	always @*
	begin
		if (rb_rollback_strand2)
			program_counter2_nxt = rb_rollback_pc2;
		else if (!icache_hit || !cache_request_ff[2])	
			program_counter2_nxt = program_counter2_ff;
		else
			program_counter2_nxt = program_counter2_ff + 32'd4;
	end

	always @*
	begin
		if (rb_rollback_strand3)
			program_counter3_nxt = rb_rollback_pc3;
		else if (!icache_hit || !cache_request_ff[3])	
			program_counter3_nxt = program_counter3_ff;
		else
			program_counter3_nxt = program_counter3_ff + 32'd4;
	end

	always @(posedge clk)
	begin
		program_counter0_ff <= #1 program_counter0_nxt;
		program_counter1_ff <= #1 program_counter1_nxt;
		program_counter2_ff <= #1 program_counter2_nxt;
		program_counter3_ff <= #1 program_counter3_nxt;
		cache_request_ff <= #1 cache_request_nxt;
		instruction_cache_wait_ff <= #1 instruction_cache_wait_nxt;
	end

	// This shouldn't happen in our simulations normally.  Since it can be hard
	// to detect, check it explicitly.
	assertion #("thread was rolled back to address 0") a(.clk(clk),
		.test(rb_rollback_strand0 && rb_rollback_pc0 == 0));
endmodule
