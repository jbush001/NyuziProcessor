module verilator_tb;
	initial
	begin
		$display("Hello World\n");
		$finish;
	end
endmodule
