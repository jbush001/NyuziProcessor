module character_rom(
	input[9:0] code_i,
	output reg[7:0] line_o);

	initial
	begin
		line_o = 0;
	end

	always @*
	begin
		case (code_i)
			11'd321: line_o = 8'd48;
			11'd322: line_o = 8'd24;
			11'd323: line_o = 8'd12;
			11'd324: line_o = 8'd12;
			11'd325: line_o = 8'd12;
			11'd326: line_o = 8'd24;
			11'd327: line_o = 8'd48;
			11'd329: line_o = 8'd24;
			11'd330: line_o = 8'd48;
			11'd331: line_o = 8'd96;
			11'd332: line_o = 8'd96;
			11'd333: line_o = 8'd96;
			11'd334: line_o = 8'd48;
			11'd335: line_o = 8'd24;
			11'd373: line_o = 8'd48;
			11'd374: line_o = 8'd48;
			11'd380: line_o = 8'd48;
			11'd381: line_o = 8'd48;
			11'd382: line_o = 8'd32;
			11'd383: line_o = 8'd16;
			11'd385: line_o = 8'd124;
			11'd386: line_o = 8'd198;
			11'd387: line_o = 8'd198;
			11'd388: line_o = 8'd198;
			11'd389: line_o = 8'd198;
			11'd390: line_o = 8'd198;
			11'd391: line_o = 8'd124;
			11'd393: line_o = 8'd48;
			11'd394: line_o = 8'd56;
			11'd395: line_o = 8'd48;
			11'd396: line_o = 8'd48;
			11'd397: line_o = 8'd48;
			11'd398: line_o = 8'd48;
			11'd399: line_o = 8'd252;
			11'd401: line_o = 8'd124;
			11'd402: line_o = 8'd198;
			11'd403: line_o = 8'd192;
			11'd404: line_o = 8'd96;
			11'd405: line_o = 8'd24;
			11'd406: line_o = 8'd6;
			11'd407: line_o = 8'd254;
			11'd409: line_o = 8'd120;
			11'd410: line_o = 8'd204;
			11'd411: line_o = 8'd192;
			11'd412: line_o = 8'd120;
			11'd413: line_o = 8'd192;
			11'd414: line_o = 8'd204;
			11'd415: line_o = 8'd120;
			11'd417: line_o = 8'd96;
			11'd418: line_o = 8'd112;
			11'd419: line_o = 8'd108;
			11'd420: line_o = 8'd102;
			11'd421: line_o = 8'd254;
			11'd422: line_o = 8'd96;
			11'd423: line_o = 8'd96;
			11'd425: line_o = 8'd254;
			11'd426: line_o = 8'd6;
			11'd427: line_o = 8'd6;
			11'd428: line_o = 8'd124;
			11'd429: line_o = 8'd192;
			11'd430: line_o = 8'd198;
			11'd431: line_o = 8'd124;
			11'd433: line_o = 8'd124;
			11'd434: line_o = 8'd198;
			11'd435: line_o = 8'd6;
			11'd436: line_o = 8'd126;
			11'd437: line_o = 8'd198;
			11'd438: line_o = 8'd198;
			11'd439: line_o = 8'd124;
			11'd441: line_o = 8'd254;
			11'd442: line_o = 8'd192;
			11'd443: line_o = 8'd96;
			11'd444: line_o = 8'd48;
			11'd445: line_o = 8'd24;
			11'd446: line_o = 8'd24;
			11'd447: line_o = 8'd24;
			11'd449: line_o = 8'd124;
			11'd450: line_o = 8'd198;
			11'd451: line_o = 8'd198;
			11'd452: line_o = 8'd124;
			11'd453: line_o = 8'd198;
			11'd454: line_o = 8'd198;
			11'd455: line_o = 8'd124;
			11'd457: line_o = 8'd124;
			11'd458: line_o = 8'd198;
			11'd459: line_o = 8'd198;
			11'd460: line_o = 8'd252;
			11'd461: line_o = 8'd192;
			11'd462: line_o = 8'd198;
			11'd463: line_o = 8'd124;
			11'd521: line_o = 8'd56;
			11'd522: line_o = 8'd124;
			11'd523: line_o = 8'd198;
			11'd524: line_o = 8'd198;
			11'd525: line_o = 8'd254;
			11'd526: line_o = 8'd198;
			11'd527: line_o = 8'd198;
			11'd529: line_o = 8'd126;
			11'd530: line_o = 8'd198;
			11'd531: line_o = 8'd198;
			11'd532: line_o = 8'd126;
			11'd533: line_o = 8'd198;
			11'd534: line_o = 8'd198;
			11'd535: line_o = 8'd126;
			11'd537: line_o = 8'd124;
			11'd538: line_o = 8'd198;
			11'd539: line_o = 8'd6;
			11'd540: line_o = 8'd6;
			11'd541: line_o = 8'd6;
			11'd542: line_o = 8'd198;
			11'd543: line_o = 8'd124;
			11'd545: line_o = 8'd126;
			11'd546: line_o = 8'd198;
			11'd547: line_o = 8'd198;
			11'd548: line_o = 8'd198;
			11'd549: line_o = 8'd198;
			11'd550: line_o = 8'd198;
			11'd551: line_o = 8'd126;
			11'd553: line_o = 8'd254;
			11'd554: line_o = 8'd6;
			11'd555: line_o = 8'd6;
			11'd556: line_o = 8'd62;
			11'd557: line_o = 8'd6;
			11'd558: line_o = 8'd6;
			11'd559: line_o = 8'd254;
			11'd561: line_o = 8'd254;
			11'd562: line_o = 8'd6;
			11'd563: line_o = 8'd6;
			11'd564: line_o = 8'd30;
			11'd565: line_o = 8'd6;
			11'd566: line_o = 8'd6;
			11'd567: line_o = 8'd6;
			11'd569: line_o = 8'd124;
			11'd570: line_o = 8'd198;
			11'd571: line_o = 8'd6;
			11'd572: line_o = 8'd230;
			11'd573: line_o = 8'd198;
			11'd574: line_o = 8'd198;
			11'd575: line_o = 8'd124;
			11'd577: line_o = 8'd198;
			11'd578: line_o = 8'd198;
			11'd579: line_o = 8'd198;
			11'd580: line_o = 8'd254;
			11'd581: line_o = 8'd198;
			11'd582: line_o = 8'd198;
			11'd583: line_o = 8'd198;
			11'd585: line_o = 8'd254;
			11'd586: line_o = 8'd24;
			11'd587: line_o = 8'd24;
			11'd588: line_o = 8'd24;
			11'd589: line_o = 8'd24;
			11'd590: line_o = 8'd24;
			11'd591: line_o = 8'd254;
			11'd593: line_o = 8'd252;
			11'd594: line_o = 8'd48;
			11'd595: line_o = 8'd48;
			11'd596: line_o = 8'd48;
			11'd597: line_o = 8'd54;
			11'd598: line_o = 8'd54;
			11'd599: line_o = 8'd28;
			11'd601: line_o = 8'd198;
			11'd602: line_o = 8'd102;
			11'd603: line_o = 8'd54;
			11'd604: line_o = 8'd30;
			11'd605: line_o = 8'd54;
			11'd606: line_o = 8'd102;
			11'd607: line_o = 8'd198;
			11'd609: line_o = 8'd6;
			11'd610: line_o = 8'd6;
			11'd611: line_o = 8'd6;
			11'd612: line_o = 8'd6;
			11'd613: line_o = 8'd6;
			11'd614: line_o = 8'd6;
			11'd615: line_o = 8'd254;
			11'd617: line_o = 8'd198;
			11'd618: line_o = 8'd238;
			11'd619: line_o = 8'd254;
			11'd620: line_o = 8'd214;
			11'd621: line_o = 8'd198;
			11'd622: line_o = 8'd198;
			11'd623: line_o = 8'd198;
			11'd625: line_o = 8'd198;
			11'd626: line_o = 8'd206;
			11'd627: line_o = 8'd222;
			11'd628: line_o = 8'd254;
			11'd629: line_o = 8'd246;
			11'd630: line_o = 8'd230;
			11'd631: line_o = 8'd198;
			11'd633: line_o = 8'd124;
			11'd634: line_o = 8'd198;
			11'd635: line_o = 8'd198;
			11'd636: line_o = 8'd198;
			11'd637: line_o = 8'd198;
			11'd638: line_o = 8'd198;
			11'd639: line_o = 8'd124;
			11'd641: line_o = 8'd126;
			11'd642: line_o = 8'd198;
			11'd643: line_o = 8'd198;
			11'd644: line_o = 8'd126;
			11'd645: line_o = 8'd6;
			11'd646: line_o = 8'd6;
			11'd647: line_o = 8'd6;
			11'd649: line_o = 8'd124;
			11'd650: line_o = 8'd198;
			11'd651: line_o = 8'd198;
			11'd652: line_o = 8'd198;
			11'd653: line_o = 8'd198;
			11'd654: line_o = 8'd102;
			11'd655: line_o = 8'd156;
			11'd657: line_o = 8'd62;
			11'd658: line_o = 8'd102;
			11'd659: line_o = 8'd102;
			11'd660: line_o = 8'd62;
			11'd661: line_o = 8'd54;
			11'd662: line_o = 8'd102;
			11'd663: line_o = 8'd198;
			11'd665: line_o = 8'd124;
			11'd666: line_o = 8'd198;
			11'd667: line_o = 8'd6;
			11'd668: line_o = 8'd124;
			11'd669: line_o = 8'd192;
			11'd670: line_o = 8'd198;
			11'd671: line_o = 8'd62;
			11'd673: line_o = 8'd254;
			11'd674: line_o = 8'd24;
			11'd675: line_o = 8'd24;
			11'd676: line_o = 8'd24;
			11'd677: line_o = 8'd24;
			11'd678: line_o = 8'd24;
			11'd679: line_o = 8'd24;
			11'd681: line_o = 8'd198;
			11'd682: line_o = 8'd198;
			11'd683: line_o = 8'd198;
			11'd684: line_o = 8'd198;
			11'd685: line_o = 8'd198;
			11'd686: line_o = 8'd198;
			11'd687: line_o = 8'd124;
			11'd689: line_o = 8'd198;
			11'd690: line_o = 8'd198;
			11'd691: line_o = 8'd198;
			11'd692: line_o = 8'd198;
			11'd693: line_o = 8'd108;
			11'd694: line_o = 8'd56;
			11'd695: line_o = 8'd16;
			11'd697: line_o = 8'd198;
			11'd698: line_o = 8'd198;
			11'd699: line_o = 8'd198;
			11'd700: line_o = 8'd214;
			11'd701: line_o = 8'd254;
			11'd702: line_o = 8'd238;
			11'd703: line_o = 8'd198;
			11'd705: line_o = 8'd198;
			11'd706: line_o = 8'd198;
			11'd707: line_o = 8'd108;
			11'd708: line_o = 8'd56;
			11'd709: line_o = 8'd108;
			11'd710: line_o = 8'd198;
			11'd711: line_o = 8'd198;
			11'd713: line_o = 8'd204;
			11'd714: line_o = 8'd204;
			11'd715: line_o = 8'd204;
			11'd716: line_o = 8'd120;
			11'd717: line_o = 8'd48;
			11'd718: line_o = 8'd48;
			11'd719: line_o = 8'd48;
			11'd721: line_o = 8'd254;
			11'd722: line_o = 8'd192;
			11'd723: line_o = 8'd96;
			11'd724: line_o = 8'd48;
			11'd725: line_o = 8'd24;
			11'd726: line_o = 8'd12;
			11'd727: line_o = 8'd254;
			default: line_o = 0;
		endcase
	end
endmodule
